`timescale 1ns/1ns
module int_weight1_bram (
    input wire clk,
    input wire [9:0] addr,
    output reg [511:0] data
);

reg [511:0] mem[0:783];

initial begin
    mem[0] = 512'h005bffba00180037ff84ffe2ffb8ffc5ffd500d600c4ffc3ffdbff61003effb60068ff47001b009e0076ff95007eff11ffdeff87006d0000fff50015004fff80;
    mem[1] = 512'hffbaff74ff62ff46003b000b00520073ff40002800d20023ffa1ffc70046ff3affc2ffecff5a0043ff780010004b004a00340079fff00015009000e3ffc6000f;
    mem[2] = 512'h000fffef007400130012007300d7003600d4ffc0ffe4000b0021ffb10046ffa6ffce00880055004f00590022ffc80054ff5d00290000ffdbffbdffea000d003c;
    mem[3] = 512'h0002002e0017ff900060006dffe5ffb1ffc500400008ff87ff2f0034ff72ff9500870096006cffd5ffe200c4ff250025005affe0ffef00a4ffee006cff8cffc1;
    mem[4] = 512'h004effdbfffa00630019ffcaffe80043ff74ffcdff930025ffb00014ff94002d0007ffce00040055ff9b0083ffd80064ff83ff83fffdffebfff8001fff64ffe8;
    mem[5] = 512'h005aff7c004900000040ffcc004d0091ff5fffe300ca0040ff21ffccff7f004e000e0018ff92ffb2001bff47ffb5007c0090ffa6003c003f004300500045ffef;
    mem[6] = 512'hfff8ffcdffb800c3007c003eff7c002aff65ffe1ff4e0039ff98ffa0003dff2e002dffe9fff8005eff5d0013002200b7ffd1ffcb0061000fffe40016ffa7ffca;
    mem[7] = 512'h000bff4900010069ffc8ffe1ff7fffe5ffd7000affa7ffb40019001c001fff3f004cffa80012005affa0ffb900bd002f0024ffc2009bff8c0024ffed00840033;
    mem[8] = 512'hffc7004e002ffff40041005f0008003bfed5ff870048ff970038001ffffaff7dffcaffb5ff30fffaffffffbc001b0027ff400091ffe4ffbbff68ff500045ff9c;
    mem[9] = 512'h00320011fff70075feed007cff570021fff3004cffc5ffb7ffa2ff40ff8dff80ffa8ffd8ffbcff81ff86005fffecff40ffedffbb006f0061ffcf00330098006d;
    mem[10] = 512'h0039ff2effc0ffb6001fffd3ff90ff49ffad0013ffbd00b6ff60fff60059fff10035ff79001a00450072ffe9006e00480088009100cfffdcff96ffbb000d0042;
    mem[11] = 512'h0027ffcd00250020008b003eff7f0069ffe2003dff8eff9c0033ff4fff97ffbd005eff79ffd90074ff5d0025002a0080002fff5200520011ffd6ffaa00300070;
    mem[12] = 512'hffcd0018fff2ffd50029ff64001100d10027006effe0ff88ffe600460093ffb10045005e0034000effe8ffebffb2ffe200e2ffc8ff6affa3004f007400080066;
    mem[13] = 512'h0047ff8900f5004a004dffb4ff89ffbaff710068ff4a007d004fffc5ffe10040006a002bffedffe50011ffcafff5fff3ffbeffc2001f0037ff88000eff97ffd1;
    mem[14] = 512'hff3bff3dffd2ff9700e9000effefffdc0018fff1fff6ff68001e0003008b006700eeffe4ffb2ffbdffe300a4002000aaffeefffa007dffc9ffc2ffabffff0018;
    mem[15] = 512'hffe4ffef00630027ffb8ffd6008bff80ff950050ffb1ff8afff6ffa6000bfffe0051ff3e00490043ffa1ff82001cffcaffb4ffaeffcd001d00eaffa8ff840024;
    mem[16] = 512'h0033ffbcfeeeff49002500100099000fff8a0057009a00d40031ffe9ff68ffe9ffe50058ffb500460091fffeff50ffe2005cfee60014ffc4ffbbffc9ffb50082;
    mem[17] = 512'h0070fffdffc5ff9affcfffb4ffe40003ff89fff3ff56ff7bffc0006eff60002400f1ff81004fff73ffc3ff270055ffd4ff7b00a7ffe7ff64ff81005affff004f;
    mem[18] = 512'h003affa0ff3f002d0093fff7000400c4ff44008000b20092ff94fffa0006ffbd002e0052ff580156ffc200300049000e0009ffdfffc8ff4e0017ffbbffcdffe1;
    mem[19] = 512'h0033ff4f005700660017002f006e0025ffd5ffb1fff1003dffdbff650007003aff98004100240096ffed0053002400d6000b004f007300df0021ffedff83002b;
    mem[20] = 512'hffda008d00daff69ff68009bffdc004d00280060ff92ffe3000cffc0ff5effb4ffc6ff330051005c0080ffa3ff9d000f001e000dff8f0045ff6affa3fff6ff8f;
    mem[21] = 512'hffe4ffda00da00350015ff41ffdeff96ff61005200160020001dfff900660126009d0064001400a30022ff59008affb5fff6007aff5d007a008cfff4ff3e001d;
    mem[22] = 512'h000efffcffa9fff9ffef0078ffbeff50000cffb00019ff76ff87ffb60120ffaeff22ffe80074ff6d00100029ffedffc3005300960062ffb6ffc3002aff79fffc;
    mem[23] = 512'h002fffe20046ffdb006100c6ff75ffa300030007ff6e003f0049ff8600eeffa500c2001affdeffa40001ffbefffc002efffcfff00000003f0077000cffeefff6;
    mem[24] = 512'h00570048ff65ffc7ff7800130039fffe000cffd9001ffffe003f0010ff54000000270031ff5eff7c00260009000a0025001fffa10020001f0030002c00520009;
    mem[25] = 512'h000dff6aff97004a002bfff0001500e8002c004b0078ffd7ff2aff60ff220071006efffaffddffcc004b0060002e000700b9ffdd00e10079007fffff00450080;
    mem[26] = 512'h0049ff9a00700041ffd3ffdd007effe6ffaeffb2ffc9ff7d00520020ffc9ff31ffbffff100c600600062fef7ff1bffbcffe20045000affcc008c000900d6ffed;
    mem[27] = 512'h0012005cffa9ff7000b8000e005e0035ffcf0032ffceff08ff30006d0018ff88ffdd0036fff0ff5800230086ff940039ffefff9fffcaff8c0099ffe5ff71fffb;
    mem[28] = 512'hffb7ffa3ffc20004007aff920086001400650044ffb9ffd9ff79ffe4000f00390005ffc000380014ffc8ffc4ffdfffb3ff81ff75ffc5007efff3001c0064ff9d;
    mem[29] = 512'hff7d00c6ffd9ffb0ffcaffb7003fffd4ffca009cfff6ff240058fff90032002800feffd5fffa0062ff9e00c5ffe9ffd30028ffb1005c006f000800d6003cfff7;
    mem[30] = 512'hff9c000eff9dfffa011fffaf0076ff93ff89ffe6ff99ffd6008fffd10039ff79003cffd8002500bcffca00250008004b002500a50097ffa900a1ffffff48fff7;
    mem[31] = 512'h009effb2000800900056ffd9ff6b007c00130048000600b2fff000370022016500d0ffdb0084ff76ffaf0029003f00750032fffaff8a003f00bfffcc003b0086;
    mem[32] = 512'hffa0ffdc0032ff60ffc7ffff001200800043ffceffc2fffd0020ffe2ffcd006dff7a00350056ff9100280017fff20016ffa9002cffb5ffcbffe4ffb0002e003d;
    mem[33] = 512'hffd1ff53ffa400280037ffc1ff9cff29007f00590057ffddff99ff9e00390090ffbaff7bffe2ff5fffa9001f00f4004a002b003bffbdffa5fff20076ff59ff1a;
    mem[34] = 512'h00030014ffd4000dffcaffc2003affbcffa8ff1d001400a1006e012dffcefff800220054ffe50086ff47ffc0ffaaffb6ffbb00960058ffed003d00b0003dfff0;
    mem[35] = 512'h0090ff68fff3005effef0044ffbc0044ffe6ff47ff930014ffd0fff60009ff6dff5dff2bffb1ff40ffab003a00350032ffec00b40018ff96fffdffedffde00af;
    mem[36] = 512'hff85008e0040ff9c00120017ff58ffd9ff2fff9bfff9002bffd0ffe1fee8005bffb6ffaa0047ffd2ffb3001600110029003900440033fff0ff64ff47ff90004a;
    mem[37] = 512'h00430046ff4100aeffc5ffa2ffd5000fffd4ffedff9400450023ffaa002c005100530024000e0020002a004cffc000080033ffc8ffdf008f0006ffdf0070ff76;
    mem[38] = 512'h004effc70018ffb800cc00430064008dffb100af006b001900af008effb300d3ffe7004fff9f003700050021005f003affabffd1ff36ffcc008c0026006b006b;
    mem[39] = 512'hfff1002ffff3ff7d0035004400140064003500470027ffe400ad0007ffdaffc6008a005fffd8ff70ffab004c0012ffb5ffccffb30000ffe1ffe800420071ffe6;
    mem[40] = 512'hffe80026000c0021ff9e0011007dffb5ffa50059ffecffdfffab0061fff30088ff2b003e00230019ffefffd3ffd5ffd5ff6cff740054ffd7fff4009e000affaf;
    mem[41] = 512'h000bffc8ffecffc90017fef40097ffad00780018ffd5ff71ffd0ff87000cff8700210079ffa5ff7aff82ff38fff6ffafff260018ff4dff7e0030000afffa0067;
    mem[42] = 512'hffc9002fffe500a6ff9500030008004fffccfff9ff610064ffe7ffc10002004e002f0055fff0000c0024003000d80028ffdcffbbff88ffcdff7f00a80070ff92;
    mem[43] = 512'h005b00c5ffc9ffe600ad002cffe50065006800ca0032fff9ffeb0038004bffd2002fff83ffafffd20047ffd40056ff70ffcffff1ffdfff85001aff08ffeb00bb;
    mem[44] = 512'h0016ff94ffb9ffd9001c0026ff6700630097ffccfff1ffa6ffcb0062ff44ffe7ff9a00e2ffd60054005bffc0ff5cff6a007dff4effb20036ff780053ff8effed;
    mem[45] = 512'h0016fff900100004fffaff76ffca00090040002f0040ffab0014ffadffe4001a0087ff7f002afff2ffffffefffd90105004e008d0003ffdd000b006fffb6004f;
    mem[46] = 512'hffcd000e001e00490003ffce002d004aff7c0021ff7dffc70064ffb0ff3f00320038ffc1ffd400ef002cfff9ffd5008500080038ffee00b0ff91ffcaff9b00ac;
    mem[47] = 512'hffc5ff41ff7fff9dffef004700090098ffbd002afff60024ffd9ffb4004d00a2ffc8ffa9ffee00acffcc00dbfff00124ffe6ffbcff61ff37ffd2ffed00440025;
    mem[48] = 512'h0009ffe9ffd0ffd3ffa1004afff3fff6ffc3ff60ffddffc100330047fff100010093ffc1001700b6ff3e008d0031006b002c0060ffe5ffe5005aff8dffa0fff1;
    mem[49] = 512'hffe0ff3bffb10006ff4ffff2ffc700020053ffa80023008e003a0037ff5700e600740076ffe9000d0046ffc4010d000affe0ffe10054ffcb0021ff9d00190037;
    mem[50] = 512'hffd50010fff1fff000960067ffebffb7003cff1bff5f005a0014ff6affe1ffc400adff7b002400180083ffbdff6eff91ffe800b5000dffd5ff9c008e004aff90;
    mem[51] = 512'h002fff68ff650054007e00080000ff70ffa70039007f006c0043009dff85ff910018002cfff7003b0059fff500b00026006aff8a00220049ffd2ffe10025ff50;
    mem[52] = 512'h00d0ffe5ff86fff2ffcfff5c00b600390048007600630009fffe0002002c006bff70ff2fff7effa1fff70045ff30004dffa60066ff800044ffedff88ffb30059;
    mem[53] = 512'hffd60015003b007d008fffa5ffccff8dff2800d9ffe700beff8c0086ff940088ffaaffd40018ff9900b1ffb4ffd70021004eff8c0007ff610060004bffcdffac;
    mem[54] = 512'hffd9ff97ffecffbfffd6ff5e00a8ff4e000c000c009800210013003b00600057ffcfffd0fff3004d00800011004afffa00510016ffc200690028002effccffd7;
    mem[55] = 512'hfff1ff4dffcb0076003dfff4ff7dff7c00590034ffc0ff7800410036ffe20023ffd50066ffcb004b0067001a00750065ffa80026fffcffbe00a300a20091ff7a;
    mem[56] = 512'h0035ffc20023007bfffb004200530049ff63003eff64ff90ffdbffd9ffd000a6fffe00be0019ff5e001200690016ffe7ff8e00a9ffa2ffd7ff42fff9ffe00041;
    mem[57] = 512'h005000b9ffcc0067ff81ffffffc00099fff7ff6d000e003c0082ffb4005bff12ffa9ffcb00770044ffcfffc8000200370037003eff26003800acffeaffe1ff6d;
    mem[58] = 512'hffdeff280057007100c500030097ffe3ffe90072ffb4fffc004dffae000600540051001eff76ffaa0041ffbe000b000bffabffbb0001ff3dff970042008c001f;
    mem[59] = 512'h002effeaffd0003fffb80031ffc5ffe5ff9dffdcff6e004c0032000dfff4ff3a00220066ff64ff1f000e00900066011dff22ff1ffff7ffc00052ff9b0091ff81;
    mem[60] = 512'hffca0090fff60015ffbf0072fff4ffe4ffcbff6400a50009fff2004affd3ffd9ffd70051ffc2ff940013ff890095ffae0069fffdffb6fff200200130ffcd0070;
    mem[61] = 512'hffaf00040010005d00ac006bff73ffd4ffb0ffcf0066004c00faff8d006b0078ff51ffe2002d0007ffd50033ffeb00390053feb80036ffcbfff0ffcd00730032;
    mem[62] = 512'h00240002ff15ffaaffcfffb10034ffdbffc0ffdfff0b007f0012ffdb0050fff0ff95000eff250098007c001d0010ff1cffabff470011ff590014fffb0007ff54;
    mem[63] = 512'h0049fffd0042ff8cff80ff61ffc1ff41ffda001b0064ffe7ffe6ff8900dbffef0065001a004dff9fffc4004aff82ffb2008e003eff530093008e004aff360027;
    mem[64] = 512'h0011ff79ffe90039ffd70063ff9eff91ffc7ffb30050001600850051004e0064008a004b011d0038fffc004600660031003e001800470024ff6eff2fffce0005;
    mem[65] = 512'hfff80046ffa9ffd4fffcffa8007bffc10035ffddfffcffbdffc2ffafffc9005d00140040ffad004c0001ffea0056005d0014ff5f006f003b00090057ffb10137;
    mem[66] = 512'h00340086fffe00580024ffa5ffcdff5e0015ff2d005100a6004b0035ff4b005900000033ff5effa3ffb9004f0036ff38004fff850067004b0005ff9bff4d0074;
    mem[67] = 512'h000dffba0048ff5a00080096ffc10004002c00800060fff0fffb0085ffd7ffc7ff85ff86ffceffbbffc0ffd8ffc80013000f000affa3ffb8ffe6ff9d005c008f;
    mem[68] = 512'h00350065ff7dfff2ffe1ffe8002f008ffff0ffd50057009effb400c5003afff100140081002effba0086fff40085ff62002eff830073001e000900bfff430034;
    mem[69] = 512'hffecffa6ffaffff6004b0063ffe20035ffec008efff700f4ff4affdfffd7000d003affb6007f0011ffe6005a002fff9c0008ffca005a001a007800a100990058;
    mem[70] = 512'hfff90060fffbffc0007d0064005e0007ffbd004cffddff5effc4ffffffc0ffc1ffd8fff9006700090062ff7800950006ff2dffc9ffe4ffe0fff20040003dff97;
    mem[71] = 512'h0062ffc6ffc400110041ffae00cd0073ffac00a7003b010fffbcffcbff89004f0033001affd0ff6900240041ffcbffc500740020ff940050ffb2ffa5ffa0002e;
    mem[72] = 512'h00750001ffee0046ffce001affd1ff2cff5100120002ffd80057004c0023002900130043005effddffeaffe3ffa80054ffd90026ff60ffcefff6ffdaffe4ffe1;
    mem[73] = 512'hff95ffb500af0084ffac007d0077ff38ff820039ff67ff8bffd50010ffe30022ffe8ffcb00c0ffafffb4fffdffcd00a8fffcff53ffdc000700b2ffd60056ff90;
    mem[74] = 512'hffe8ffc7003effbe0043ffe1fff8fff30079ff3a005dff870013ff2e0041ff1a001fffed0053ff15ffe4006e00310019ffacffed001000030020ffe7ff60fff5;
    mem[75] = 512'h002dffd9ffc5ff5fff74004bffe8ffb40015ffe9ff63fff5002a00590021fffdffc90009ffcb002e0020004d007c0099ffe9ff82007cff44ffec00c10015ff4d;
    mem[76] = 512'h008cffbd001500defff40096ff7bffa4ff6fffccffa8001f0001007700040067009fffd600ab00a700160066009cffc8004000c8ff63ff2affc6004f0007003a;
    mem[77] = 512'hff99000a0019002dfff0ff750053ffe000760018ffe1ffce000bffc400450019004000ee0025ffd3ffe8006bffe30002000fff82fef0ff7b0024ffbdff4e004a;
    mem[78] = 512'h00aeffc3ffb5ff7e0042003affd800ae00770016fffbff88008ffffb00430061fff6ff85ff4cfff2fff9ffecff8fffdb0021ffb8ff0a000300920041ff3e0068;
    mem[79] = 512'h0039ffb5002c00500028002dffc9fff2ffcc00030005005000c2ff75004c00300019ff8effd4ffe500520069ffe8fffe00130021ffae0061fff0ffa1004e006d;
    mem[80] = 512'h0074ffa3005900a5ff98ffd40017ffcd0061001cffb100400029ff89ffe0fffd001700730016ffac003affa8ff95fff6ffaaff96000900780042ff82ff8b0020;
    mem[81] = 512'hffdc008e0033ff85003eff2dfff3003300900082003e001eff8dff30ffd10027ff9b0032ffbaff3a00710050ffe9004a0031ffbd0012ffa7ff94ff3cffbd0012;
    mem[82] = 512'h00550070009000810021ffdeffe4002affb200230054ff8fffb9ffdfffa8ffff001f0069fff800620015ffb7fff3fff0ff9cffb4ff78ffe20051ffb5005fffc9;
    mem[83] = 512'hffc5002400670000008c006f001d008b0094ffdd000fff84ffc80022ffc0fffffff4ff0a0023ffcc003cffd7ffbf002effdb000c003cff8affecffd9006c0013;
    mem[84] = 512'h003e003bfff2ffcfffd5ff05003c0095ff4fffcbff0a005100460073ffc9fffa0013fff50032ff7affdf0034ffbaffda00400086ff4effff0031ffe5ffd20000;
    mem[85] = 512'hff64ffeeff98ff74ff70ff95ff70000e0030001100980026000b002f0021006aff8c002dffdd0025ffca0040ffcdffcbff1f0040ffb5ffac0036005e0004002f;
    mem[86] = 512'h0014ff770044ffbbffd2ffdc000300460029004aff7a004400af0045fff900260056fff500420045ffafffd1001fffc100a10012ffc6008d000c006800800030;
    mem[87] = 512'hffbfffd7000b0019ff98001f004dffc4ff9c007d00220061ffacff49006800040042fff1ff09ff7b004e00390062ffba007000690058000c000600860027ffc7;
    mem[88] = 512'h001800610083fff7ffdc0025ff95008affdb004b0019ffb9003800d3ff6effba0036ff850043ffd4ff650012ff4a001c0131fffb003bff8effedfff7ffeaffc6;
    mem[89] = 512'h008b0082ffac00810006004500600018ffa5001b000300400022006effe7003f001eff66ffc50055007100a3003c00b5fee0ffdb001f0039004affc8fff2ffb4;
    mem[90] = 512'hffb200150076002fffd300a4ffa5ffb1002c0059ffe5ffdb00440121ff8affd8006800520013ffbbffc4ffb80019ffa70011ff9affee001600b5ffa8ff89001b;
    mem[91] = 512'h0040ffb50057ffb1003200110060008300fdffed002fffc1001700390040ffeeffe9009affb1fffb0011ffb60094ff5800c4ffc7ffcdff680017ffa700500024;
    mem[92] = 512'hff68ff7dff8aff600092ffe40037fff30029ff7cffe2003bfff500af003c0048005bffdaffa9ff830022009bffd70065ffbd0056ffe8ffc7ff9c00acffd900b3;
    mem[93] = 512'hff680057001bffbe004bffaa000300310047004900f8ff97fffdff73ffc600190075ffa60008ffacff7fffe4ff770067000fff40007700ceff8dfff7fefc006e;
    mem[94] = 512'hff60ff35ffec00a3002400530113ffdd00f900cfffcd00a5ffe4ffc1ffd7ffc0ff9100bf00840019ff96ffba002300020034ff81ffb1ffdbffb40012ffc7ff76;
    mem[95] = 512'h00490006005600e7ffe5ffb300880087000b0064ff8affeeffb1ffb4004a001fffc5ff9700bb008100cdfffc00b7ff28ffde00150042ff9effcc001f009cfffc;
    mem[96] = 512'h0028ffcfff73ff9cff9b0035ffc90078ffc60037ffa30055ffd0ff7bffbaffa9ffef009afffaffae005dffe4003bff84ffedffa4ff760005ffb7000d009bffb5;
    mem[97] = 512'h00220002ffaa000d002900250034fff60016ffb500250034ffe9ffc2ffccffdefff600b2009fffb1ffe30027ffc7fed7ff3d0055ff6a0034ffa8ffc4001f00b6;
    mem[98] = 512'hfff6ffd6ff8eff5cffc700710072003600bbffbeff48ffe7ff81ff79ffa60029ff77004aff980033001effd0006b002bff3cffffff5f0069ffe8fedc003effe0;
    mem[99] = 512'h0017ff5f0005ffeb00610066009fffe400ccffc40064ffe80023004e0061ffe6ffc1ffec008e0092ffe5001500b5ffe8ff8f005cff8a005eff290008001500d1;
    mem[100] = 512'hffd7ff3a002cff9000d3ffcc007ffffa001f00080010fff8ff540028ff94ffbaffe90083ff8cff7f00460062ffbfffc000afffa8ffbd0051ffbbff92fff5ffdb;
    mem[101] = 512'h0085ffbcffa1ffbfffdf0065ffe9000bffb10021ff7700be0014ff8b0008ffe0005e004fffde009b0023ffa80121ff5eff81003500c4ff50ff3bff5d0072ffc5;
    mem[102] = 512'h0009ffecff9200dc0052ff8c00c4009b0003006300abff96ff60fffbffcbffaeffd7ffbfffad00a1ffcdffd20116ffa6ff7afff5005cffc7009d0047ffc70003;
    mem[103] = 512'hff78ffb00036001cffe8ff47ffa3ff98001eff430069fff1ffb4000e00230089ffdf006cffd800500040001700940060ffc9ff4f00c4003dffd3ffab0080ffbc;
    mem[104] = 512'h00ae000c0003ff86008e0006fec50033ffc5ff9d001effe8ff78ffd50037ff6d0050005200f9ffcaffa7001e0027ffabff240001ff900030fff500140069007c;
    mem[105] = 512'hfffeffbaff8dfebc00a4ffb8ffa4ffec00100021ff6f00a1000affbbff46fffbff9cff890040ffb6ffc800b8001a0078ffd9ffb9ffe5fff1ffc8009affc8ffd3;
    mem[106] = 512'hffe00004ffb0001d00f6fffe006e000a0064ffc1fff6ffe0ffebffe400d20060002bfff2ffe2ffdb008b0095011fff73004400180005000fff4600800049ffa5;
    mem[107] = 512'h00060079000affa00058ffa4005bffeaff9eff55ff9a00a7ff6d00890041ffd8fff6006affd5ffb5ffb70086fffcffa9ff3c00a0006eff81ffa0ffbaffd10071;
    mem[108] = 512'hffa2ffd1ffceff7fffefff48004600590047002affd6001affc1005affe8ff890000fff00041ff09002afffe006c0050000c0006ffa60014ffbf0002ffbc001b;
    mem[109] = 512'hff330007ff92ffd8ff6200bd0030ffa2ff9a001effe50036ffdfff3e0026002fffa1ffd0009900570023006d0067ffd4ffeb00250066ffc1ff9700a1ff95ff93;
    mem[110] = 512'h0059006dff54fffaff99ff72ffeafff2fff70083ffbaffb6005effa7006100220007ffa30061ff8a006fffec00450016006bffd90014ffca001d00e4ffb1ffe2;
    mem[111] = 512'hfff20038005f0019002ffff6ffccff620098ffb6ffb0002e00a7ff7e00bfffb1fffaff67ffa7fffaff6dffc8ffffffecff72ffc3ff37ff5d00b100220059fff6;
    mem[112] = 512'h006b0078ffb2007affb3ffe1fff8ff98ffcbffc00021ffc5007a000dff68000d0074000effd10019008600330032003e00c0ff520008ffbd00ca000effa00033;
    mem[113] = 512'hfff50004ff9affbbff98ff6bfffa00bc00110060fffdffedffb9ffa3ffdaffb2ff51001700730028ffdf00920004fff4ffac0042009dff4a0094ff84ff820003;
    mem[114] = 512'h00b8ffd1000d001cff22ffe5ffc100360064ffaf0007ffe2ff8200450052ffd4feb90009fff300acfff2006a00ca0050ff72ffffffabff92002a0041ff6e0019;
    mem[115] = 512'hffc4ffea0043ffd9004affd500570101ff9d0014ffe3ffbc0017fffe00210060009f0025001affe2ff8effe0ffffffe4fff8ffe9ffad002cffe1ffe5ffcbff19;
    mem[116] = 512'h0029006e003a0058ffc1ff8000230049ffa5ff41ffc5fefefff80042ffebffdd00d5fff0ffdffff200280044004aff5c001c002cfff3ffacffc8ffd300b60006;
    mem[117] = 512'h000dffc9ffefffa8fff5ff71ffb30046ff81ff8bfff9ffe3fff6ff65ff9affbe006eff35003aff1c0018ffc7ff65fff80079ff91ff3e006c0039ffbaff87ffb2;
    mem[118] = 512'h00c5009b001000b80064ff760057ff930053ffbd001d006effc700590007ffbcffe3ffc3ffe9001bfffaff6bffde005dfff0ff0a002f008affc900a2ff9bfff8;
    mem[119] = 512'h00620001fff0ff7effe8000eff9200840008ffa40085fffb000bffbfffa9ffecff6effecff4ffffa006500650019ff680000ff42ff9b00a60069ffa3ffc0ffcb;
    mem[120] = 512'h004affe700a5ffad003affc30005007c0009fffd003cff99007affe40060ffb3001100a70014006a006b004500b40021001c0012ff3300390034001d004c0017;
    mem[121] = 512'h0029010ffffeff450017ffb9001c004bffebffdf0052ff31ff7fffdeff620074007301040014fffa0008ffda00d8005b0002001d002a000400ffffa400070021;
    mem[122] = 512'hff6c004b00d5ffd4ffb7002dff9cffe2ffdd002dffa6ffb4000affb3ffbb0047000a008700520084ffe9006d0044005cffdbff8dffbb002afff700850040fff1;
    mem[123] = 512'h00680094ffc6001e00c7ff83ffcc0025002e002d002bffdb007fffc2004800d4ffcc00fb014d0027002bffe20005ff07ffac0016ffdcffe200520035ff6100ce;
    mem[124] = 512'h0008ffecff28ffb30027ffcf0061ffa70055ffff0049ffe30024008600080007ffb60062fff80037ff70fff3ff82ff5400040013ff50fffeffbaffe9ffbf001c;
    mem[125] = 512'hfff1fffeffe3ff5eff65ff91ff78fff40016ffaeff70ff93004500110050003800ab008f0030ffcbffe9003effde000d003bffaeffc60042fff5ff57ff56ff78;
    mem[126] = 512'hffd80053ffa2005effb00071004400900006ffcfffbbff49ffe6ff7cffc8ff74000b0033ff68ffc6ffa100310049ffe5ffec008aff600056ffd2003b000bffde;
    mem[127] = 512'hff9f001aff7cfffc0045004fffae0006ffe500ae007fffea0043009eff55ff760077008dff99ffbbffe5009d0135ffd4fff20013fff60009ff95ff1fff31003b;
    mem[128] = 512'h002200ebff2e0058ffabff96006500a2ffd1ff87003700a90042ff8b002fff83002e0008ff89ff8a0009ffe5003affcf0009003fffb70005ff9c002e006effcc;
    mem[129] = 512'h00100022ffcb0021ff9e006e0008fff3000e0070005fffc2ffcb006800b30089009cffefffc30002ff9d0086007d0037ff8f0010007affa20036ffe6000c0021;
    mem[130] = 512'hffa900190024fff800a900c90025ffe7ff5b00760049ff380003007e005d0023007500bbff990035ffb0ffd5fffd006a0046ffd60009ffc60040ff9fffa8ff5b;
    mem[131] = 512'h0016ff70ff7b002fffd1ffd5fff700c4ff60ffad001ffff7ff9c0086feff0055ffedffe100050087ff800013003b0095ffceffd300100008fff0ff8aff56ff97;
    mem[132] = 512'hff90ff99ffc1ff5600dc00a00010ff8cff760003ffdaffa5ffbc0041ff910042ff4affad00b1ffdaffc9ffb3005eff7affdffff2ffd7005c001c002cfff0ffd9;
    mem[133] = 512'hffc50018ffde006900200117ffacff74ffab00310017ffa90019ff76fff10023ff5dff9d002a007e0067ffd6ffbd0074009b009f004effab0022ffb800680025;
    mem[134] = 512'h0005ffb100530072007c00620023ffccfff900b80014ffdeffa40069ffcdff63ff9bffe600160029ff92006800e8ff5afffe00420080ff8b00610048ff8fff90;
    mem[135] = 512'hff840074001a0066002f0083ffc60088ffa1ff450068ffe3fff7000f0063ff7d0058fff0ffa0ffbf00bc001f002dffdc0005001fff8cffbc007500b40055ffaa;
    mem[136] = 512'hffb70069ff9a004c00530055ffc9001aff81ff75ffbe002c005affc6008effdaffb4ffd7fffcff93004b005300510012ff91003800bbfff900abff63fff6ff8f;
    mem[137] = 512'h003effc8001fff9fff95ff8a003affec001aff89008cffd70056ff30ffbaffdc0053ffaf009cffeefffdffdf0016ff3cffe50039003bfffc00550018000d0023;
    mem[138] = 512'h005900a4ffeb00d7ffd1008d0051001bffbc006300b60017ffdf00150018ffb6ffff0044ff91007b00570007008500240008ff5cffc90034ff3700630002ffdc;
    mem[139] = 512'hffefff87ff37000c0019ffd8ffeb005c00120003fff600950044ffd200540010009800dcff6dfed1000c00a2ff500084ffb0ff60ffadfffc001b0049ff88ff8c;
    mem[140] = 512'h0027ff9f0013ffbeffd10021fff70081ffe7ffa7000bff5e0051002afff2ff850047ffc0ffc300210008ff90ff9affeffff0003fffe2fedfff7eff9bff8cffee;
    mem[141] = 512'hff08ffda00400045fff200680021ff37003bfffe000fff12008efff40070ff79ff0a007000b7ffbdffd8ff9dff93fffb00000030004bff970007ff600046ffec;
    mem[142] = 512'hffabffdbff79ffdd0074fff8ffca007cffffffe4000afff8ffaa001300180056005e0019ffbd006a0044ff5bff6a006b0083fff2ffadfff80009ffda0042ffbc;
    mem[143] = 512'h0060ff91ffb3ff5a00fdff76004fff9eff4400190000fff5004f006effe10039ffae0036ff7200b4ffbffff3ff9f003dffe200600015ffdb009200600080fff5;
    mem[144] = 512'hffdc007cff9b003cffd80042005aff65003d0083ffbc0016ff8bff960071ffaaff7a005b00f4ffc6006a0047ffbd00100008ffe1ff71008bfff0005efffeff4e;
    mem[145] = 512'h00b8ffe90004ffb8fffdfff5fff9ff69ffc1fff60092002f00750065ff8800540040000bffe3ff8ffff80093ffceffd800a0004c007100610077002d001d0059;
    mem[146] = 512'hffecffcc002fff75ff87fff7ffd3000800e50012ff830036ff3fff93ff9800500083fff0ffa3000bffbdffc5007effe2ffb70027fffe0028ff8affcc00b00098;
    mem[147] = 512'h0070ffafffb3001e008c000affef00c90039ffb7ff5eff9fffb60008ffeeff980035ffa4ffbb004a004a00570046005a0000ff5bffbb001c003700350005005c;
    mem[148] = 512'hfffb0066ff63002a0090fef7fff9004eff14004effce001d0009ff8c0058ff97ff590043005dffbfffb4fffeffe9004000440002003f0032fffdfff4ffe9ff83;
    mem[149] = 512'h002d003a002b00410000ffd5006000450043ffb4005a0082ffb9ff31ff21001700510079ff8fffe0ff7a007affd4ff9dffe6ffb6ffa60036ffeaffddffe1007b;
    mem[150] = 512'h000b000effc0ff3aff76ffd1000200b6ffeb0085001bff6e003e005dff42ff97ff8e013a0067005d00320085001aff8700e8ff95000eff6a006affa0001f003b;
    mem[151] = 512'h005f0050ffdeffb4ffd1ffa70005fffd00000012ffe5fff2004d007effeb00760023012400ddffaffff0ffe00069005300c7fffa004e0091fff60031002bffa2;
    mem[152] = 512'h005c0003009200a8ff9f0057ffb30061ff74ff30000dff7dff8eff3afff4ffb7008c003bfff8005dff6fff63ffa000b2ff8a0046fffdffc7001d00d3ffe7fff5;
    mem[153] = 512'h0015003c002d0015ffc1ffbeffb9009dff9f003fffecffccffcaffefffd900290098ffb1ffe9003f008c002d005dff31fff7ffc2001cffe00093ffa3002f006d;
    mem[154] = 512'h008cff950021002b006fff8cff4300a6ff3aff5e00b6ff34fff4ffcc0008ffb000630051005c005c000a00320054ffebffc5005b0065007fff7700baff7b0043;
    mem[155] = 512'h00280045ffd70003ff3dfff7ffbf0007ffc7ff7c006dfff200efff3d0061006700890059ff8e0038ffa50032ffeb0026ff5cffd3ffa6ffe4ffbf006100e5fff3;
    mem[156] = 512'hffc100e6fffe000400c900380001005c0060009fff4fffb2fffe001400660046002c007c00a100680029ffd800d7ff520029ff440051fff2ff7f0077fff3011b;
    mem[157] = 512'h0046001dffd6ffb9ffddffd6ffb100d7ffb10027ff7effb2ffec00c2ff2afeee002e001aff9cfff5006e001500ceffeeffdd003c00acffc9ffd000ab001c00b3;
    mem[158] = 512'h0064000c00230043005200f4ffe8001effffffddff46ffcbff69007200330098fff4ff4e0029fff4002b0093005affa7000dffb9ff920045ff340029009400ea;
    mem[159] = 512'hffca00d5ff93ff3bffb0ff0d0049ffb200460040ff9601170067ff2effbdfff7009c009b000700650001ff3400470080fff90007ffff000e007400a1ffe90083;
    mem[160] = 512'h007a0062006b000aff46ffa2ffd80070ffe200d2ff8effd8ff9c00740055ff8d0086ffc0fff7fffdffe5002300bf001c0002003e007a00b0ffb30049ff80007e;
    mem[161] = 512'hfff7003d00890033000a00b3ff7dffd6ffd20056007bff97000effbb0021002d004500caffe5ffebffb000ba000cffd80008001fffe20009ffc5001a00470024;
    mem[162] = 512'h0057ff6f00ce0019ffcd005dffc80040ffad0054fff6ffe400170069ff8cffd9ffc40075ff40ffb9000dff8b0022fff1ff97006b013dfffbff9c00d4ffcd0021;
    mem[163] = 512'h002cffc10005ffecff5400370007ff110075007c00430006002dffcb0060ff1c000bfff2ff5dffc5002e0004ffa0ff9bff99ff78002effaffefeff8eff27ff4f;
    mem[164] = 512'hfeee005aff9a004400dd0041ff800011fee200e5ff670041ffdcffd1ff8d002d0036ffedffb9ff89ff86003a00570038006effde008600dbfff8ffd5ff880078;
    mem[165] = 512'h0015ff94fffeff830106005a00150000ff4aff63ffd200e7ffdaffe1ffdc00450039ff6b0007ff4cffd8ffeaffc8000c0041ff950095ffd60053ff7afff60047;
    mem[166] = 512'h005800530004ff5eff96ffe7ff9c007cffdafff3ff6d0038ff0cff770088ffacff7d0014ffc0fff9ffd2009dff86ff9cff9700200077006e0074ffaafff700bf;
    mem[167] = 512'h000aff8effe6000dffc0003f0044ff9e00f5001dffe50048ffd8ffa2fffd0044ffb80037ff8d001400c200a100a4000dfec9ffd7001b004b0008ffea00070027;
    mem[168] = 512'hfff300020050fffaffd6ffc2ff56007bfff10044000affc3009eff8aff3cffb2ff81ffe50044000aff6effcd0055ffcf001c006200c40027003d001e0054ff66;
    mem[169] = 512'hff86002fffd000520068ffb300a8001b00370061003a000d0013ffe2ffba0080ff8affd800bf008e00a1ffa8ff94002bffacffd8ffe2ff7cffd6ff9000220021;
    mem[170] = 512'h007efff80072ff23fff90057ffde001b0003000a000fff4aff6700260000ff9f0044ffff0075001300f00009ff83ff6a00b0fffdffed0061ffd3000d0075000f;
    mem[171] = 512'hffb70006fff7002affa6008c00650076ffdafff1ff98006affb0003affb0ffe10081ffc5fffeffea00010091003f0033fff1008eff9f012c002d0083ffd70009;
    mem[172] = 512'hffccffd7ffa0ff9e0059ffefff91fff9ff9bff5dff1e004c004e000f0090006dff940043ffbb007dffca0068ff34000d008dffa8ffd4fffb00caff7f0010ffa4;
    mem[173] = 512'hfff4ff95ff49ff5e006eff9f00010090ffdcffe9ffba001f002b0086ff540057ffffffe0ffe3001f005effde006d000500670013ffff002dffc7ffb100620033;
    mem[174] = 512'h007b0024ff82ff73ff61001a0040ff23ffeb0002ffb4ffa30049ffe5ff940070ffe80001ffc6ffc4006aff950084007affab0061003cffc30080ffe00073ff75;
    mem[175] = 512'h004affdc006effaffffd0009ffc6007b002800240029000d007000410005ff91003b0026ff91008a0096ff7d00690048ffdc00250055004b0015ffa30021ffd3;
    mem[176] = 512'hff5d0017ff4e0004ffe9ffbdffee00170024ffca005f00100154007aff3d000cfff9ffab0031ffd1ffce0034ffdeffb000edff4f0015ff64ffccff8300870037;
    mem[177] = 512'hffa2ffe1ffc10048ffa9ffe4005e00b0ff96ff7bff7a0055012e003fffc7ff850009ffbefffdffba00080117fffd0054ffbe001700a8ffc90049ff8600aaff69;
    mem[178] = 512'hff5000190081000b0072ff71002a0038ffc7ffde00200022fff7ff9500970047006eff79ff64ff88ff890020ff200040ffd3ff720060ffaaff48ffac005000c6;
    mem[179] = 512'h007500790024002dfff0ffacff970098ffc7003dffdeffef00a4002e0020007e0057ffc500b30027ffc7007a002cfffe001b0062ffdcff7f004a0011ff9eff5e;
    mem[180] = 512'h002ffff90071ffa6ff9d0011ff8500740012004e0070ff5000d2ffca00b2002f0010003cffeeff9fff3500600037ff81ff890037ffe600e3ff8effb8ff97ffb5;
    mem[181] = 512'h00fd004cffbc008300400031ffd800650024ff720029ffb6fff700d7ff61005cff660036ff9a005dffadff7cffb4ff6efff500850034ffc7001f0003ff89fff2;
    mem[182] = 512'h00a8ffcaffe70095ffa50033ff290080fff3002efff1ffcf00180038009d0083004ffff7ffaeffbbffe20011004700c1003c001dffe6004600c6ff3600430004;
    mem[183] = 512'hffa40023ffe7ffd60020ffd0ffcf00c0ff8e00170050ffbb005900a50116fffa000b0044ff94ff7cff49ff720032ffd2fffe00a7005fff52008a0001ffe0ff59;
    mem[184] = 512'h0000ff55ffb1005effb20056ff7f002dff6b000c0020feb90029ffd6009efffcff85001e00370022fff7ffffffe20008ffbd006b00adff4700b5ffec00520040;
    mem[185] = 512'h0076003fff9efff200040066ffec00b800560061ffe3ff69ffd90026006d0066ffd1009afffbffdd00aa000fff50fff30093005bffa9fffdff4bffa6000ffff4;
    mem[186] = 512'hffc800b1fff4003b004b0009ffe1005a000eff9f0065ff60ff99002f00220022fff600350096ffe90063005a002c000f0030fffbffb6feb201010038ffe3ffce;
    mem[187] = 512'h002b0016003d00310071ffc6ffdf00bd007a0039fff3006d004ffffaffbcfff3fff3005800890031004e0079ff53ff6b003cffe9ffe8ffffffac007dfff60020;
    mem[188] = 512'h00b50028007c002dff7c00ccff7d0006ff8d001e000dff46ff2300a4ff6fffadffc3ffa3000000380029fffcffefff6affc600abffffffaafffbffe9fffa0030;
    mem[189] = 512'hffa80087ffa0ff8affb5ffcbffba002700370094ffe20026ffe90016ffaa0029ffa90065fff1fff4001bffbb00c30023ff9fff91ff69ffde004700310020fff5;
    mem[190] = 512'h001600150049ff38ffeefffcffb60078ffc60010ff660083ffd1006affe8ff870038ffe6ffed0023ffdd00cb000c002e002b001d00560059ffeb002700300004;
    mem[191] = 512'hff9afff1ffecff9aff99009affe2ffb1ffbdfff6ff960096fffc003c0003fff1ffcefed0ffe4ff9900e20017003aff90003f0022ffcd00a9fff0ff88ffccffbc;
    mem[192] = 512'hffa7007effad00e9ff580010fff200c600000038ffd6000e000c002d000affcc004100d40068ffdc00170044ffedfec100300063ffecffefff8700450007ffc6;
    mem[193] = 512'hffcaffa5003bff53ffc7ffbd0043007aff37ff58ff9eff3fffcf0026004a004e00630102002cff95ff41ffbb001fff980092ffee0010ffe7003aff95001fffd3;
    mem[194] = 512'h003d002d0079ff44ffeeffccff8e003affb40018ffb3ffedffbe00390084ffa0002dff4bfffd007dff090012ff2c0052001dffde00d600c0001f0061002e0027;
    mem[195] = 512'h00a6ffee00310007fffc00bfff1b006cffffff79ffdaffb70014ffc30017ff980001ff5bff3f0003ff9a00500094001f0025ffa7ffbf0090ffb30015ffddff7d;
    mem[196] = 512'hffe6ff96007cffc2ffbd00300048ff9affa0ff8eff1b0064ffb900410022ffddffa7ffa30011fff800730011ffcafff4ff84ff7100530025ffd8ffb3ff7200ad;
    mem[197] = 512'hffa4ff9afff2009000140028ff83ffa8ff670018007400280014fffaffde00a80004ffc6002eff8b0025003aff5bffae00160027ff82ffdefff9ffd1ff9c002d;
    mem[198] = 512'hff2c004d001fff64003d00530057ffc90098fff5ffdeff52ff9fffeeffc6ffac0057ff94ff42ffc20010004200070050001fff9affceff9fffb9002a006500fd;
    mem[199] = 512'h001dff9b0100ffcfffcd0027fff000150074fffbffd50058ff99009100df001cfff3ffe6000e0075001b00be0066002aff9a00070039ff6dffbf00b90012ffad;
    mem[200] = 512'hffffffd50016ffd800b5ffc0000c006affdf00620054fff5ffa2002cff4b0063001ffffbffe8003e004dffb30018000d003fffa0ff75001bff6e0002ffd5ffd1;
    mem[201] = 512'h000cfff8ffd60048ffcaff930020ff8d0053ffd8004cff40ff85ffe9ff8f0069ff1e008afff9007900790065000f002c0032ffd80022ffeeff50ffc000ac0005;
    mem[202] = 512'h000b001a00470035fef500070054ff940020ffd2ffe8ff6bffec0056004400190047ffd7ffa9008600bf000d001900210065ff36004affbbff7c0032000aff7b;
    mem[203] = 512'h005bffe400160067ffdd001500a3009b00420016ff6afff000b2002400060033ff7d006fffe0ffdeff9a0025001efffeffd20068ff6f0024ffb3ff99ffccffa2;
    mem[204] = 512'hffc70021001fffecffd3ffabffa3ff600025ff8b008e0072ffb1ffa3ff98000cffaa002500efffa00012ff950044ffdaff3dff2e0030ff95ff26ff750069ffd6;
    mem[205] = 512'hfffbfee3fff10054ff3cffc5001c00daff9e0026ffef0002002f003e001900290050002b00130003002400280047004e003b007affb5000e008b005500fa0055;
    mem[206] = 512'hffff0067ffc8ff38ff3cff910052ff8cff68fffeff5eff53005800340059fff20028009f004d000800690020001effd9ffa8ffd6ffe2ff3e0010ff9f002d0019;
    mem[207] = 512'h0006ffc5ffb20020ff49ff94ff390018ff9cffd9000d0058ffe000e700960077ff23001f0014ffb20072ffa40077ff95ff90ff0a001dffdcfff1ffc00002001c;
    mem[208] = 512'hffc7013800560006ffda0077fff30091ffb5fff10065003c002f0077005800830024ffe5ff72ff7dff29002a0018003fff9bffa9003effa5006c0001ff8bff30;
    mem[209] = 512'h00040001ff6200fb0059ff27ff9d009400160003ffa8ffc80031007300f2008cffc6005800850002ffd3ff720005ffd8ffe1ffe1001b010500a7ff4000330054;
    mem[210] = 512'h0023005600020032000a0046000d0025005a0031fffbffc2007a0021008300b500300063ffa7fffeff3cffefffab00d2ff820099ff97ff3cff34ff8a002200a1;
    mem[211] = 512'hfffa006cff9fffad0054ffd0fffcfff4ffce0023005affe4ff82008801100037ff9600470000ff8f00fcffa50064000effea00060068ffebffd4ff3300730071;
    mem[212] = 512'h0023006cfff8ffcd009dff95ff2fffd1ffd400da007100820097003a00a8006dff770016fffd00210037003cff33004cff72ffaeffd60006ff82ff7f000affbc;
    mem[213] = 512'h004cfffcffc3ffbfffdd0027002b004cff570074002700b6005800b700cf007afffb00c5003900aa006dfff6ffd8001e0047ffb30025ff5c0005ffe2005dfff5;
    mem[214] = 512'h0084ffd0003eff6bffbcffce004900fe0043005e0094ffa9ffe900cb00ddff89ffad0006fffffff9ffff001a00170002003b00a50069ffae01040022001a007e;
    mem[215] = 512'h002bffd3ffc1003effc20074ffd8009effa4ffa4003b00acff91008c003c004e000c0048000f00580096ff74ffc40029ffdc007affd60037ffffffa5010bff9f;
    mem[216] = 512'hfff70080ffc3ffc4009000b3001e0093ff85003c00e10039fff1ffef0039ff74006bff04ffb300bc002dffd400c800a20075ffd600dcfff10065004affd7000e;
    mem[217] = 512'h0012007fff050107ffc6ffb70091ffc900550077ffbaff78007400d00096ff95fff1ffc4ffcbffd3ffa4fff6ff7b006b002000460032006e0062ff9affc1ffeb;
    mem[218] = 512'hffff0000ffc4ffb10012ffadff8b00ac0014003affbbff670003ffd0001affa7ffb5000b00320082ff75ffac0009ffa2008300420049fffa0086007cfff30022;
    mem[219] = 512'h002a001c004bffaafff00086ff9e0062ffee0049005600980082ffc7ffb00017fffb006a00270046ff9e00a2ffcfffda0014fff5005cff9a009700a8ff85ffc7;
    mem[220] = 512'hffdaffb7ff73ff93ff59002800cafffa00140033ffa40007003d009dffd8002d0016ffab00660039003b006400eeffe90066000100a9ffc10030fff0ffc6ffe3;
    mem[221] = 512'h001e0055ffa6ffbeffe90053ff6000030030ff70ff7f0038ffb9ffb7ff49ffd200dd0027ffc6ffa2ff6600740052ff6e003000120012ffbc006effba004eff85;
    mem[222] = 512'h0003ff75004fffedffa5ff90006300340050ffe4ff48ffe3000b0057ff62ffbaffb3006cff02ffd0002affd4ffe30071ff8eff7f00330014000cffbcffd100cb;
    mem[223] = 512'h001f004e003c0028ff57ffd7ff90001d000cfff3ff98005f000eff6a00170026ff2b006a004b0044ff77003200660014ffe7ff93004fffedffde0071fff2ffec;
    mem[224] = 512'h00700012001400d2003b0011ffc7ffbe01030001ff71000aff600097fff7fffd0090ffefff39007e000a00190004ffe2ff4d001fffb0ff4dffad0056ffb1ffff;
    mem[225] = 512'hffa5ffb3ffaeff74ffedffc50006ffed006a00a10081feb3009affd9001ffff0ffcf00800021ffeefffe0025003dffd2000dffc4fff5ff1cffb7ff4b00510096;
    mem[226] = 512'h0032ffe3000fffe20031fffaffdcffea0070000f001d0025ffc5001400cbff72000effff001e005aff98005fffef0039ff49003a002dff40ffca0068ff9fffb2;
    mem[227] = 512'h00c00031ff9c001d0064004e002000740043003bffcc0011ff3b001200230049003e0046ffd500c6002dffc80038ffe300390002ffb4ffcb002e002b0014ff40;
    mem[228] = 512'h002aff9fff9cff91ffc50019ffc3ffc80021ff82001fffb6ffac00350059ff400003ffa5ffa600cdff880082ff73007affbeffbdffdbffb8ffe400260071ff2f;
    mem[229] = 512'h00c8fff5ffe300040066ffe2ffa60005000d006e0047fff9003700170098003e0093ff9a006b00050029ffbf0031ffa2ffe700b6ffdf0025003200dbffc2ffa3;
    mem[230] = 512'hffd4ffa8001d00420003ffe8003cff3aff82001a00040011ffdcffe60042009200a0fff700bcffeafffc00180005ff86ffbe0051005a0042008c006a00abffea;
    mem[231] = 512'hff870074002dffc5ffc6ff96ffc00020ffc5ffaeff750066004dff7cffa4ffc4ffde0026ffbeffde007eff74ffa800e800a4007dffbbff1affdbff9a006a002a;
    mem[232] = 512'h00850006fff3fffe001bffc70003003a0022002900390021008c0083004d0056ffbcfffbffccff5d0033ff57ff96ffc2ffffffe60069ffea005f009effa7ff3d;
    mem[233] = 512'h0099ffefffc7ffee000dffb3fff4006e0042004dffcefffefff300c9ff8a0028ff82001b00d700210031011b0066ffb1ffb5004b004400900063ffed0088ffe3;
    mem[234] = 512'hff450004ffbaff76ffacff920058002aff9a00ab0002fffbffa4ffeb000a008d0061002fffabffd00015ff50ff5c0017ff9f002effebffdeffe40056ff7c0013;
    mem[235] = 512'h00400084ffdc001bfffa00870058ffccff6b000ffffeff72ffc1012600a40004001f006c0082008bffdfff8300a1ffa1ff50ffe100240019005900490034004c;
    mem[236] = 512'h009affed0069ffaa001eff56008000090083ff9cff21ff9c007600ccffcb0043ffe8ffb8ff6bffe7005bffe100420040ffa7007f0022001c005affdc008a0041;
    mem[237] = 512'hffdf000f00410020002e005d00590078004ffffdffed0046ffeeffd200890073004affd4000effc9ffbbff82ff97000fff730001ff8d0050000b0034004e0059;
    mem[238] = 512'h00cc0029fffcffe5005500450048ffee003cffd8008effd9ff7f006f003c00ee00860024001400500056ff50ffc1006c002a0079ffd2ffc5ff38ffc1fff0ffa5;
    mem[239] = 512'h0050007bff6f00b5ff8fff78ff1a0055002cfff8ffc8002e0094001f008800b1fffb007cffe0ff80006f001bff37005eff6c003dffe0ff450006ff910037ffbd;
    mem[240] = 512'h00360088ffe1ff9200330050001f00900013ffb700e300840018005100ab0063ffb40042006800a7ff75ffb0ffa5ffa1fff10006000fff7f000a007fffe5009a;
    mem[241] = 512'hffb00005fff3ffe2ff33ff61ff37ffb1fff1011b003a010500290009fff3001cffff0043ffed005201050050001f0046ff8300edffe400770039005d008200bb;
    mem[242] = 512'h002ffffcff50003a0018ffc70010ffd50022007f0143000c000b0029009a0072ffb90015ffadffe10092fff6ff64ffea0024ff4f0054ffe60011ffb6ffe7fff2;
    mem[243] = 512'hffa500ea00dffff40004ffd3ff81ffac00af009d00920062009ffff9ffd5ff6bff2d00a2ff880075ff74ffba001600a300e1fffeff8e006cffe10090ff87ff8c;
    mem[244] = 512'h008bfff4008cff8bff83fffd001100af003f004b0089007f004dfff6ff970021ff35002efff4ffa50029007affbf0061ffeeffcbffdc009700a1ff6affe7ffc0;
    mem[245] = 512'hffbc0015ffca004bffa90049ffca0029ffb8005800aa008f0048ffd7ffcf000afff3002b00600005ff98ff880054001aff9bffea006dff7cffaaffc9000c0073;
    mem[246] = 512'hffda0000ff930067ff9bfff8fffd00ad00340085ffaf0077005cff96ff6aff3fff5e0067fff9ffa9ffbdff8cffc700870041ffc50046001b0071ffb000000087;
    mem[247] = 512'hffb700bd0027ffefffb00039ffb5fff200690028ffe6003dff91003fffca002b00d4ff4300cbffccffcf0066ff90ffb3ffe5ffc5007e00dcff8dfffb006c005b;
    mem[248] = 512'h0001002a0069ff9dfff8008c005f00b20049ff5600b5ff8d00780067ffb2ffebffbd0037ff85002effe9ff97003aff96005000c9fff5003c0014fefdff7e0046;
    mem[249] = 512'hffe0ffc700d1ffc4ffd1ff5f0018003c0053ffd300850064ff58008affec00a2fef70024000affb6ffb7ffd2ffff002800070047000fffe90072ff94ff820089;
    mem[250] = 512'hffd3ffe00011002dffea00370019ffec0015fffc009bffbbffc1001a003effa3ffe1ffec00200033ffe0ffe1ffae0040002600080053003200c1007dffbe00bb;
    mem[251] = 512'h00320035ffbdfffcffd4ff50ffc50031ffe9ff9dffe000290040ffe9ff3dffcfff1000b1003c0047ffb50005ff9a008900400024ff68ffa3ffb800520076008f;
    mem[252] = 512'h006000310045ffc1ffd5ffd2000eff82ffd3003f0070fefe002a0019fff00071ffc6ff7fff98ff7dff81ffa6ffc9005e006f004e0096ffcc009effc50076ffc6;
    mem[253] = 512'hffe4fff100beff3e001400040003ffda001fffb2ff8cfff400650032ffa0002dff64ffe3002cff35ffe00033002f0008ffb70018009effd3005cffc20008fff3;
    mem[254] = 512'hfff50096000cff640028003bffdcffc5ffbcfff7ffce002affd0003cffe7ffedfffa0063001d0023ffedffdc0043ff50ffdcffdbffc8001a001000c7ff82000b;
    mem[255] = 512'hff53ff6a0010ff99fff5ff52000bfff9ffcf00080073ff510044fff20064ff800066ffce001a0013ffc10022ff6f0078ff9f0016ffbd00a1ff7fffaa003d005d;
    mem[256] = 512'h00bc0039ffd6ffd10055ff930055001600120051001e005bffd0ffe9ff94ffdeffb000ebff5dffe1ffdeffe5003f00240032ffaa00350007005dffb4ffe2ff56;
    mem[257] = 512'h005effc8ffd0fff1000bff9eff5e00a40041ff6bff94ff7fff510005003700090067fff7002dffa100ff003f0028008cff28ffa1004fff0cff01ffe1ffecffde;
    mem[258] = 512'hffb9ff6d003cffa6ff8bff8e009a00eeffa1ffe9ffdbff2d00580052ffcb0058ffd800240007004b0010000d0025001bff1c005900010050ffde005b00590066;
    mem[259] = 512'hff9e0068ffe5003efff3ffbdffbafff9002c0001ff6d0082005c0006ff3e005b0072ffbdffec0025ff580053ffd3005500490080001e00250024002dffa00035;
    mem[260] = 512'h0028ffdbffe00065003cfffc0071ffd7003800670020ffb000640028ffb1ff9e00c3ffdc004f0009ffb8ffa1008900760011ffa70049ff3500eeffa80032006a;
    mem[261] = 512'hff97001cff1a004dffc9ffee008fffadffc2ffc5ffacffdb00510065004d003c0068000401340001fffb003bffe10110001600e5ff8f00b1ff940045002ffff3;
    mem[262] = 512'hffbfff30002b001e00a5007d007dffab003200af0034ffef00b40070009e0036ff4affd70021ff140058ffd5ff9f0026ffe0002900e9ffaaffdf00a700760091;
    mem[263] = 512'h005bfea7005bff94ffadfff6010c0111ff4c0037ff51ffd80023ffde00780034fffdffb8ffaaffc10083ffdc00680073ffcfffe70002005dffc0002a0026ff98;
    mem[264] = 512'hffdcffc10045ffdfff9fffcd008b0060009f00480023ffdeff17003a004f006effa500820029003a00710095ff210095ffdbffe8001bffab00abff8500240099;
    mem[265] = 512'h0000ffcaff8d006a0031ffcf006f0038ffb900ca003f008b001e00240029003e0053ff5101140047ff620040003aff9effd9000300a3003d007c007e00420009;
    mem[266] = 512'h000600d1000900170002000d0081002dfff3ffe1009d00c400a40030ffc2007a006000d50017ff98001dff9dff9d0060ff520036ffcfffa100b30035ffb2ffe6;
    mem[267] = 512'h0028fff6ffc8ffc9ffe70015007c00450027ffe3009affffffdc0069ffdf00560041007c00c0ffb90040fffb0032ffd20000ff22ff6ffefeff68ff92003dffee;
    mem[268] = 512'h00c1ff3effc80024004b0027004efffe00b4ff79006600d900bc00beffadffce00e3003fffcdff8b00b90013002f0041007cff89ffffff95ffd4ffb200940042;
    mem[269] = 512'h00070071ffa200efffb2ffe4003200380076000700ab000affe0ffe8ffc7ffb300720083ffd4ffda006d000fffdd0052ffa9fedaffdcff93ffa4005cff65ff9f;
    mem[270] = 512'h001f00aeffd700a4ff8bffe300440067ff82ff8dffe6004f008d0077001fffc400550042ff5bffa90068008bffca0020ffb5fffdffd3003c004400c6ff850067;
    mem[271] = 512'h000f0051000000c8fef5ff3fff9a007c0077ff5400460101008cffb60070ffc7ff7d00150062004500720017fff9001dffb6002b000700880071ff9effce00c8;
    mem[272] = 512'h002d00bd000d0043ff78ff84ffdd00220013ffe100160086001fffcfffb9ffda00bb003d00370061ffabff81007b0072ffef0031004eff4fffe500c8010700a7;
    mem[273] = 512'hffb30023007d0066ffafff51ffdbfff9fffc0040005efff400a4001500250073ffd1000c00480081fff200bc007affc80065001aff9e003b005affdaffc20072;
    mem[274] = 512'h00270050003e000fff9e0027ffca007a00caff78003e00890001ffd8fff90077005bffd7000e0009ffb3ff66ffcb0029ffe600210001002700720036009b0023;
    mem[275] = 512'hffb8fff5005bffe3ffc900010030ffc70073000f0045fffefffa005cffae000a009fffaffefc002d004dffd1ffd4ff2fff7200f6ffe5ff330098ffe300240090;
    mem[276] = 512'hffceff4a00e2ff91ffe8fffa004f00840051009eff770017000e0000ff1e0007ffacff70ffeb00c1001bffafff38ff9500460036ffd300b7ffc4ffea00430002;
    mem[277] = 512'hff95ff930017ffc9ff68ff3d00a2ffe8ffedffdf006cffacff89ffe0002dfff80039ffc7ff9aff6effed001200a2ff97003900a7ffa7ffe3ff4dffb10025ffc0;
    mem[278] = 512'h008cffad004100010014ffd400f50031ffa4ff7b005a0007004c001cff530022ffe5002e002b006a0089ffd3ffabffbaff96ffb50003004cff9efffeffe2ff53;
    mem[279] = 512'hffedffddff97ff87ff4affcd005cff620091ffb1000f008affad00a60064003cffd8ffd2000c000dff6e0020ff7e0064ff77ff18002cfff3006dffe2ffe7ffab;
    mem[280] = 512'hffdcffdc00baffd60018fffdffb4ffa70069001dfed50086ff95ffa100cc0070ffff006bffdc004400eaffd5ff390025ff4300270031ff62ffb500b9ffcbffd6;
    mem[281] = 512'h000f002d0020ff09ffa5ff89005b0011ffd1ffe8fff40039008f000cffa2ff7fffe000680023fffcffa7ff70005d0033ff47ff3600bdff78004dffccffe70059;
    mem[282] = 512'h00280025fef400baff6fffa20013ffb400b7ff61fff7ff5500130020005bff130087008a0001fffffff300a8fefc00e90084002fff34ffea00100066fff4ff03;
    mem[283] = 512'h001e005500880010005affdcff8c008f00390018ff85ffd7004eff60002b000c002affeeffac0030006f0078ffe9003eff420037ff4400150052003d004c0043;
    mem[284] = 512'h004c0085ff960074fff20057ffa2fffaffe600a90002ff7b0002ffffffceff6e000f0066ffd400350068005d0037ffa1ffcd0008ffa2ffb2ffe300040045fff4;
    mem[285] = 512'h0024ffb3ffc60025ff18ff0f00c6fff2fff3ff5effe2ff9d00050079003a0034001eff550046005aff810028004a000bffd80029ffdbff5bfff8002700960014;
    mem[286] = 512'hfffa00530058002400380069ffe5ffddffd200cb003affff005100960020ffdb0123ffe600cdffe900c2ff980015fff1003d007f0067ff9f0007ffe5001eff84;
    mem[287] = 512'h0002ff660044fffcff8c000d0052009eff86ffb7fff3ff4afff6003a00810039ffa6fed3008fff92ffc1ff88ff6a0046ffa1ff85006c0003ffd2000d0015004e;
    mem[288] = 512'hff33ffa1005200270036ffdc0033ff9f00b60040ffb7ff59001aff8a0020ffd80058ff3d0032001e0002000d0003ffadff69ffac000600b40007000a005c004d;
    mem[289] = 512'h002dff4b006c000cffa5ffec004000940085001cffc0ff85ff46ffd0ff9e00390008ff4000abff9a000c00a0ffaaff8effc1ffaa004900870071000effe2ffe1;
    mem[290] = 512'hffbe001a0024ffd200d10024000a0067ff6000e2ff83ffc000890080006600550068ff19003100080061002cffc2007eff65ffc800bcffe8014300ad003effb2;
    mem[291] = 512'hff71ffb10058006400340094000affe2004fffeaffc0ffbc00590018fff5ff68ff7dff33ffdfffed002f0004ffe60008ffc0ffd9003900060066ffff0031ffee;
    mem[292] = 512'h0007000bffe4fffeffea001b0079ffe00085002dff8bffd400290092ffb6ffaa0025febfff83ffdbff7bff89ff83001aff990088fffa00ff0034008aff94ffd8;
    mem[293] = 512'hffec0003ffb50010ffcdff67ffffffa8002effb5003c004d002d0032ffcafff6004aff7dffea003a0064ffee001b000d001300b900160017ffc2ff9000130052;
    mem[294] = 512'h001b00440095ff7d0063002affeefffd008bff9f005b004d0027ffdeffb90035fff1ff38ff660021ff8bffea0020000aff46004400410085fff0ffd7ffa1ff75;
    mem[295] = 512'hfffc0073ffc7ff9c003dff9f00eeffc8ffd8ffad00a7013a00820053ff650086ffaeff9a0069002500e500930071ff7eff73ff67ffd3ff6a002b006c0043ff94;
    mem[296] = 512'h001c0076ffe50007ff1700410147000a0011ffe300cc0005fff0003b003700a1fffd00dafffe0003001a005f004d00c10036fff5001c003b0029ffa0ff67ff98;
    mem[297] = 512'h000c0000003bffbbff610048ffd800220046feb7fff6006bffb00009005b005c0014ffec002fffc8001cffc3ffd200b4ffc0ffca00640059000a008300defef6;
    mem[298] = 512'h00a8ffd70056ffad0025ffb1fff4ffad0058ff83007d000a00a900f2fff50003ffec0070ffd6002700a9ffbb0027ffae0048ffca0080002effadffb1002d0034;
    mem[299] = 512'h005e00a700240088ffd4ffe6ffc0ff50ffbb002500350049ff92000f004d0074ffbd0022ffb6ff7c0000ffb4ff99005dffc6000fff7a00530025002d0013000c;
    mem[300] = 512'hffc8fffa007c0053ffceff64002cfff1005aff8100adffbd004c0086ffccffa5ffefffe5fff00008ff240024ff6a0016ffcb001300b8ffe70018000affd500dd;
    mem[301] = 512'hfffaff9cff7f0046fee3ffc500b00008ffd7ffcd010600760083ffb7ffe10068fffb00bbffd200caffdb008900390058006c009c00bfffd1005f0000ffef003a;
    mem[302] = 512'hffb5ff46ffbf00e800780062006c0072000f002effdb0074000b00040044002200d2ffdf0017ffd40042ff7cff94002e00360029003dff4e001fffe2ff86007e;
    mem[303] = 512'hff310041001d0018ffd700500074ffb50008ff93001fffc3005300d1008effc4ff8bffb000f0ffe10060ffe9ff6cffa6ff790089ffe6001dfff9ffeaffe700a2;
    mem[304] = 512'hff9affdcffba001e004a0010ff75ff900008ff51ff700092002cffbbfff70025004affd6ffa1ffd5fffd00400063ff610059ffd60029002b0034005bff83ffde;
    mem[305] = 512'h007900310052ff10ffc3ffc10061ffb0002cfffa0045ffe2ffa90062000fffaa0026ffd80026003aff7a002effca0009000d008d00070012ffb40018ffa40069;
    mem[306] = 512'hffebffb70004fff5ffe5ffe90009ffc2ffb7ffa7005bffa10041fff4005aff09004400abfffb0077ff650065ff950037003e001f0009ffda0081ffd2ffeb0040;
    mem[307] = 512'hffd800030027ff1b00690058ff8900b5ffdeff58ff2bff6dffa9006c0043003600a0ffac001b002800700029ff1d0007ffb1fff2ffc7ff9c00aa006d0063ffdf;
    mem[308] = 512'h000b003200e80089ff29ffa60016ffa9ff8700170087fffd006aff5dffaa0036001b0141001b001f005300190018ff9fff7a006e00dbffe4ffc1ff3cffd2008b;
    mem[309] = 512'h005fffc2004dff95ff5fffb5ffc50050ffad000dffd5ffdaff07ff9cff950024fffdff980030ffdc0022ffb6ff78fff1ffceff690026fecffff7ff29ff5effa4;
    mem[310] = 512'hffc0ffb6ffccffe7ffb0001c0038ff7cff98001afff100eeff910059002fffb300120071001afffc00d4ff64ff530028ff3e0095ffcaffd3ffe0002effd50034;
    mem[311] = 512'hffeeff1affb800320055ffc7ffc80067006bffef0041002f00360123004a0058ff64ffcbfff6004d0046ffdaffbfff4f003e00a70009000effaf0023ffcbff9d;
    mem[312] = 512'h0017ffaefff7ffa2ffafffc9ff84ff97ffbdff3e0099ffaa0041ffdb002e0049ffb0ff6e0057ffe3001cffcb00180044ffb00004005a000cff72ffd90087ffe9;
    mem[313] = 512'hffd9ffc5ffe2ffe7ffd4000f006c00360002ff26ffe5ff5cff99ff70003f00d6006cffb7009eff56005dffffffd6ff53ff90ffc8ff91ff4fffaf001cffc3ff97;
    mem[314] = 512'h0056ffad00750014004c0085ff2e0014ffc60007ff680031004a00de007f0008ffcdff9f000f000a00c1ffc9ffc1fff80020fff6ffc2ffa1ff59ff9800b3ff8b;
    mem[315] = 512'hff45ff37ff32ff8cffac000cffc6ff980053ffdbffaaff4600a3006000000035001dff19000e00c2005b004f002ffff3ff610070006b000f00220086001f0022;
    mem[316] = 512'hff5300190037000fffa0002a001f0030ffa6ffabff500003004d000700480055ff76ff8dffdbff1cffbcff83ff9d000b001dffa2fffaff04fff2ffe60053006d;
    mem[317] = 512'hffcc004d002000c4ffbe00acff7affeaffebffbcff6eff3f00fe0082ffdd003cffd1ff4affe6ff9eff49ffd6fff20029004a003b001b00670070ffe200570064;
    mem[318] = 512'hffeefff7ffe50089003e002effc1ffeeffb0ffc50016000dffe20055ffd6ff660054fea70022003cffa1ff4b002f003affff007a0011ff980082005e0000ffde;
    mem[319] = 512'hffc5ff5fff700090ffef000b0018ffddff5b00680075004e005fffc300540008000bff25004fffcd001d00320077ffd5ffdefffe0034ffda0017ff8fff6a00a0;
    mem[320] = 512'hffd200c5ffbe002d001b00b2005cffe1004bffeb007e00a9ffe1001f0000ffeaff6ffeea001eff8fff17ff2d002affdd006aff94fffd00c7001200f0ffa50005;
    mem[321] = 512'hffc3fff40039ff6aff830089009dffacffd3ffcd005affbaffb70022ff7e012cff91ffc1ffde0038ffe0ff99fffaff81ffd00057ffb10001ffec00560039016f;
    mem[322] = 512'h0039ffa6ffe0ff9e0014fff400a9ffdc0056ffff00990045008d00960014ffcaff89ff8afed4ff70006dff6300830035ffbbffc4ffa4001b008cffec0007ff95;
    mem[323] = 512'hff8f006effccff58ffc000b4fff0ff82fff9ff40006300abfffaffb0ffbf00a8ff63002eff3e0020fff8fffbffe2ffd7004e003ffff0003a00710042ffe80003;
    mem[324] = 512'h006dffba005bffddffb9008f0033ff9a001dff7100a6ffe2ff61ff7eff81006cff9f007affe0ff50001e005b007fffd7002bff7e0061ffc80065002c00d1ffb7;
    mem[325] = 512'hff53ff21ffaaffbbff52ffc90006ffdc000effa50039ffeeff29ffd0000c0040ffcd0015ff94ff740010004c00640089ffd5ffef00c500730049003500690065;
    mem[326] = 512'h0019002aff82006aff66ffb3006f00a0ffe1ff4000b1003200dbffdffffcfff6ff6e0029fff00047006400e3ff41001e0066ffaf00020011ffc5ff18fffa001a;
    mem[327] = 512'h00290040ff9b0008004000350010ff0cfffaff8100c9ffc40024004d00d100bdff81002a000b0029008f001e0022002400b0ff510053006a00300034002bffd5;
    mem[328] = 512'h001dffedffe200bc0080fee1ffef0007ff9afffb00240023ffc8ffff0089ffee001dffdd00580078fff6fff5ffff00dbff9b0016ff6d006900420062ffd1005f;
    mem[329] = 512'h0009008200b4002f003f00540054ffa7ffb2ff0800d9ffd00003ffe00073ffebfff1006400bc008500030017fec5008eff8effecff69009b001a002f0038000c;
    mem[330] = 512'hfffeffe4ff9d00faff840025ffebff98ffd9ff5d00320064ffbe002d0002001fffdf001f002f000c003affacffe0ff95ffc6000b00390082ff38fffaffa40072;
    mem[331] = 512'hfff80008006bffac00090090ffa00009ffd1ff460035ffed001cff9aff80ff6600a900070058005900290019003a0039ff28fffd0020ffbb0052ff9e0027ff7b;
    mem[332] = 512'hffabffc1fff700110067ff81ff49001b000c0088ffe3fffbffce001bffc3ff80ffb50040ff91003f003b0046ff5fffb6ffcfffff0008ff65ffef0053ffa4ffbe;
    mem[333] = 512'hffc6ffa4ffc60011ff44ffee00060010ff8b0041001300720024002affe2ffd6002d0083004bff1b0040009600410053ffc3004bffad007d001effc7fffb0072;
    mem[334] = 512'h002bffe100040012ffcfffe3ff71002eff58ffd10011ffb40025005d003ffffd0053ff91ff86000b00160008ffef0010fff3ffca00070003ffdefff1ffe6ff2a;
    mem[335] = 512'hffb3ffc80079ffff0000ff94000cffbd00a500a0ff6d007e008d0020ffe7006a00af0036fff00016ffa4000e0000ff960007ffb3ff90006a002b001d0005000c;
    mem[336] = 512'hffdbffd3005b004fffaeffe60029ffb60046ffec002bffc7ff6cffe0fffc002fffa8ff87003affadffe5ff5efff300790040ffd2ffea0040ffc9003fff75ffe5;
    mem[337] = 512'hffba006cfff8006effd1002effe5ffb8ffe30084ff61000cffdd00260000ffcc00420009ffb7ff3e006fffe40019ffcf0084ff77fffd00a00020001cffdaffa3;
    mem[338] = 512'h0092ff8dffc5ffb1ffd100290014009dff6affd70078fff3ff7c0014ff8fffdcffd2ff57ff7900140028fffcff9aff960071005eff9000580027ffcd00bf00a3;
    mem[339] = 512'hffed0048ffcb0048001c0003ff570002003600060045ffa8ffa9ffa9006800450028002bffc7004affc4ffc700250055fffbffe30044007800bbffc7003d0020;
    mem[340] = 512'hff810024ffa6005a0010ff93ff9bff770023ffe100660041ffbbffeeff7400b4ffebff6f000a000fffb2ffddfffdfff2ffcaffd4ffcf005a007cff2dff4d0025;
    mem[341] = 512'hff6fff6d0049ffa90030ff55fffbff98005e0037004fff89ff04ff86003aff9b006c0019006fffa10029002affdfffa5000b0027ffce0084ffdd005c00a7ffea;
    mem[342] = 512'h0017ffa60056ffc4ffc90053ffca00940033ff600068001d0007fff8001300720049ff4bff97ff9d00710017003b008a003fffe8ffd1ff92002a00a8ffa0ffe9;
    mem[343] = 512'hff4eff6effe9004e008e00010070ff750041ff75ff4b0044ffbeffc90015001cffabfedbffcb009b0072ffa7ff1fffb0ffb700d9fff0ff2f00aa00010020ffbf;
    mem[344] = 512'hff5bffb70024007fffa1008d0079ffbaff8aff6d001dfff00068ffd600e7ffc8fffeff51000a0084ffe6005b004fffe6ffebfff8012a005d0072007b007d00d7;
    mem[345] = 512'h003c003eff5cffc6ffe8ffc30043ffa0ffb1ffbc00160052001f000b00abffd2fffcff3fffbd0007fff900a7ffe9005d00ffffb60045ffc5009f0054ff76ff1e;
    mem[346] = 512'h0067fff70060002affe10091003affe100cd0001ff9a0030ff840017001a005affe6ffc0ff7400370012006e0049ff920042fffa004a0046001bffe4002efffe;
    mem[347] = 512'h006d00460050ffe4ff510039ff6c006affce009900120097ff57ff7afff800e6ff8dff6b008300170021ffc60030009700c8005d00d1ffbaffdf0035ff650018;
    mem[348] = 512'hfeb1ffca0063000b002000a500680018ffd600250003ffd6ffe5ffa50005ffc7ffc0fff3006bfff9ff9fff8b00c4ffda0084000d0063ff8ffffaffc2ff9b00c3;
    mem[349] = 512'h001a003affc5ff93ffee00670035feb2006c0009fffa0031ff4b00a5ffca00bcffe7ffa20051001effe7ff52004aff58009f005fffc4ff63007a005fff7c0071;
    mem[350] = 512'h0035ff88ffd70015ffde00f800000045ffbe00260057000100a60004003100920003ffaafeefffb5ffe90023004dff910088ffc9feff00a9fff4008c0003fff6;
    mem[351] = 512'h0094006fffa6ff6f00220099001dffdf0018ff13ffe9004a00b6ff74ffc400ff001effa50013fee90029000f0001ffef002dffdf0038fffc0089006900770033;
    mem[352] = 512'h005f000400040022000bffb1ffdaffbbffa0ff1bfffa004a0001005e004b00e00047fffd002dff8fffffff9e0046003e00d7ff8c0011ff1f00630029ff8f000e;
    mem[353] = 512'h0046fee1ff95ffb900570006ffe7ffa60031ffd50000002700e0005a0071fff80046ffbbff6efffb0002000bff9600ebff8eff9effeb00160005007200d7ff8c;
    mem[354] = 512'h00aeff71ff7d0053005affd7003fff7800b2ffd900abffb1ff520059ffc100350037ff590043000b00b1ffe30012008affa4004d000500490062ffcc00bbfff4;
    mem[355] = 512'hfff6002a0068000e0048008affeaffddffd0001a0007ff05005b00660011ff51ffe00055000cffccff87ffeeff6d009e001eff8700fd001900750015002f00c1;
    mem[356] = 512'h004dffef001400220008fff8ffe9ff56ffa7ffbb0069ffe3002600570036ffc8fff6ffe6002100110007005f001e00b4ff4eff5dff94ffcb001a006a00ad003b;
    mem[357] = 512'h0004ff7d002fff08003bff24ff2bffffff5fff64ff90ff56007dff8bffbcff9afffe00720065004c0056ffb00004fff6ffe2002cfff900ce009fffee00150049;
    mem[358] = 512'h000b005a001800bb00cf0029ff9affd100a6fe88003dfff7fff200e200c1ffff001cff7afffe0096ffab001500480083002cffa4ffdbffca00b400260021ffa9;
    mem[359] = 512'h001d009e007fffcb0027fff80021ff720005ff42002eff71fff4ff680096ff79002cff13ffc400c4ff71fff9ffc4ffffff91ffe2003c0056ff1cffc4ffb2011f;
    mem[360] = 512'hff8d00230059ffbd004bff3fffd8ffaaffc20017ff7e007afff4000700110042ffe5ffb800320077ffa7ffc3ff6dff7700a9fff20042ff24fff0ffe300820109;
    mem[361] = 512'h005fffdeffecffda008e0008001d002100520029005e00550073ff50ffd200140047007aff68001cff970057fff7ffb9ff36fff4ffc5ffeeff61001ffff00037;
    mem[362] = 512'hffdf0074ffafff8cffc3ffa70079002affd10020ffeaffdffed400b5ffba009cff870089005f002bffdd0036ff910031ff6600490003005c00260006ffdaff78;
    mem[363] = 512'h00030011ff4100040038002eff9affb7ff920021ffb8ff85ffae0030ffc6fecc004ffff801300006000c0017004b00bf0088000dffb2ffbdff98ff66ffdaff95;
    mem[364] = 512'hffb60024ffb7004300bf003cff98002000850059ffff0045007bff38004c004300e0ff9f004d0051004cffc600c1ffe7000b0002fff00086ff3affec0042ffb8;
    mem[365] = 512'hfff8fefbfff1000fffc7ffc2ffbbffe9ffedffb9ff92ffd7ffa1ffc9ffaaffa30048ffa0000b004effd60042ffd10071008fff8cfff80064ff4cffb40041fff4;
    mem[366] = 512'h0008ff65ffac005c0016ffe60069fff6005cfffeffc2ffb3ff83002dff7dff52001a003b0038ffc7fff0005500450035ffc3ff85ffb10015003b0079ffeaff6e;
    mem[367] = 512'h00a5ffd7fffeffc1ff98ffa9ffa3ffd2ffc40074007fff86fff7001100330008ffffff710032ffd3000effe9ffb5fff4ff740012ff0cffdc00300063ffa4ffcf;
    mem[368] = 512'hffd2ff70ff8c00480015ffd2fff5ff8effb30027ff85ff7a00440098ffc8ff8f008effa20087ff79ffbafefaffb0ff82006b00970044011dffe5fff00016ff90;
    mem[369] = 512'hffde003dff7800bdffcc000c004a001a00b9005400bf000effbd00320050004fffbeff7bffb40001001affaaff76009e00740048002e0023fffe003affbfff1e;
    mem[370] = 512'hffea007dffe90016fff4ffdcffbaffc0009bffa6ffe10060ffb9ffc10064ffdaffceff0300a5ffd0ffd7fff400a4006dfffcfff3009200b20014000b00350030;
    mem[371] = 512'h00350041007f001bffabffac00bb002dffb00029ffa5fff8ff69ffd8ff50007a005bfe8effe20008005fff90ff9dffeeff8700180051ff6b0005ff77ff4c003d;
    mem[372] = 512'hff920038ffeb000d0081ffecff67ffe5004d003f00280027ffb0ffbe005f00a6fff2ff5cffac003a005dffbeff6d000c002fffa500bd000c0013ff9d00caffa7;
    mem[373] = 512'h0002ff65ffa5004ffff2ff8800dd003e002600130019ffdaffc60004ff82ffb9ffa1ff2200d00044ff8f0059000400160055002fffde00c20096ffbfff930012;
    mem[374] = 512'hffa7ffe5ff43ffac0027008d0002ffca0070ffba0000003fff800024004cff66009e00100070008bffe20010ffc800150053003200b500bcff3efffcff17ffc9;
    mem[375] = 512'hff6affd6002000b7ffc200180025004c006b002bffcd0094007a00880078ffb6ff14000500a40026fffc003c0000ff7300f7ffcd003300e7009b0056fffa0069;
    mem[376] = 512'hfff4ff660111ff610015ffb400640024002e003cffeaff1d003aff990075ffc000050046ffb8ffa6ffcf0120008afffd00a9009a0073ff4dffc4fff1ff72000f;
    mem[377] = 512'h001fff3e0006ffaf00080078ffa7004fffd9003cffc80028fff6ffc90103000000280053fff50033ffd7ff85ffef0007008f0100ffd40002003d002affda00a6;
    mem[378] = 512'h00fb0050ffccffa6ffa4007100c60013ffa30032002d00160092ffdafffc006affb4fffa0040ff8fff8affe9007d003001220002fff2002400bc001300f20043;
    mem[379] = 512'h001d0065ffbd009e013f00fa004c0008fff40022ffb4ffddfffe0015ffee003d0004ff9effdfffd6fffbff8cfffc00b5006eff720006ffe6ffbe0016ffde0004;
    mem[380] = 512'hfff0ffd4ffc000c8fffa004affffffaa00020043006fffe1ffa6fffb001a0075ff87ffaafff6ffb5ffc4ffab00a40122007d0038fff2ffdc0001004f001affaa;
    mem[381] = 512'h00d7ffc0ffedffc2008300390004ffcdffd10025000b0021002bffe80077ffa4fff2006cfffd001d0023fffcff9200320150fff0fffdff8e001c00720037002b;
    mem[382] = 512'h0038ff970096ffb50056ffe8ff6b00d3ffc300290054ff94ffc4ffeb004f007bff320007008fffb5ffac00a70089005f0072ffea00390033005bff85001affa1;
    mem[383] = 512'h002600120010006dff5dffdb00a40005ffc5ffe00024ffcaff4effec005200bcffb0ffa40039ff8dffe10043002f00db00160023007000ba00500066ffca0007;
    mem[384] = 512'hffabff65008bfff4003c00a1ffacffcbff89ffe8ffe7ff78fff50097ffc600c300130013007c0090feb8ffe8ff7dffefffe4ffc600380038ff950049005e0055;
    mem[385] = 512'hffa8ffefffa300d6009000a20099fff5ffe9ff4fff4bff7effe7ffe90082004dffad003cffc200b2fffdffed00260021005cffc90031000800090032007bffd7;
    mem[386] = 512'h002900a3ffb200390028ff7eff9aff79002b000dffa0ff9cff9b0022ff9700250080005f001bfff500b0ff42ff7c004affefffc00059ff70002b001c00d50055;
    mem[387] = 512'hffde001b0025001a005effacfff1ffc5ffd7006ffff2000c0043ff9affc7ffde00e0fff500bdff5effa40004ff6effc4ffe6ffe000150098ffb5fffc0093ff7e;
    mem[388] = 512'h0043ff88002d00190012004e0021ffc7ff7c003a0061ff87ff8b00b700090044ffb4ffd70049ffe9ffe40024ff21ffeeffe5ff91009affcd00a5ffe8ffe5ffa8;
    mem[389] = 512'hffcd002effc5ffcc0056ffcdff1b00110005ffe90058000aff170033005e0008ff9e0047ff6c0000007affd2ffeaff48ffd2ffb0fff1004effd80023ffecffd3;
    mem[390] = 512'hffd1ffdffff8ffc10039001cffca005aff80001affbcffc7005d0027007cff24ffe70050ffa900490007ff40ff9b00270087005a000e00990061ffdeff47ffc5;
    mem[391] = 512'hff90ff9900810009ff8f0040ffac00a0ff48002b001dff53ffecff5b000fffcfffa6ff53ffed00200056ff7500720022ffb4001d0040ff95ff7effd20070ff58;
    mem[392] = 512'hffabff82ff8e0058ffb2ff85ff80007b0059ff89ff7aff5600bdffb7ffd20048001e00240038ffe90033003affcffff9ffbd0055fffd0043ff7300fc00210089;
    mem[393] = 512'h0041001d0085ff56ff37003c0055ffb4ff1bfff5ffdd00b4ffe80036ff51001afefdffa5001effe4ffbfff7dfff400860065ffeaff8affd4fffdffee00f0ff51;
    mem[394] = 512'h004effed0092007d00500084fffb0044fffdff5bff93ffd3000b0060ff68ff4e002dffc2000c003fffe3003e0016ffe2008d00420020002cff73000f0001ffb6;
    mem[395] = 512'hffa3ff770027ffd2fffc00390022002a001300e3000bffdfffd6ffa4fff5ffc2ff77ffe5002f0010ffd3ffd7fff400eb0048ffc5ffa7001e0017006b0049ffda;
    mem[396] = 512'h006f0067ffb10098ff940008ffb5000b002900090006ffbfffb5ff8aff33ffd800020032ff9b002bffaa001d00a1001c002affa8004cff5700e30003ff8bff77;
    mem[397] = 512'hff9dffe0009d000d003dffaf003fff960010ffd3ff8c0033ff8aff8effdaffe60073ff5effc000540040ffbdff6b0036007f007e001900310008ff77ff61001e;
    mem[398] = 512'h000dffe70084006affb20028fee4ff74ffd8ff58ff65ffdeffe6001effffffc8ffb20096003fffbeffaa0161ffc1ff8000c7ffb4004dffeaff650007004c0079;
    mem[399] = 512'hffbc000f0092005f002c003fffc2ff93ffdb0009ff9cffd40020005200adffc8ffe3ff54ffb90052ff50001dffd2ffb70024ffd1006bffd500360063ff76ff81;
    mem[400] = 512'h00e1ffb0ffd000150081ff53ffe7002800f40046ff41ff35ffa1ffe80030005fff74ff930036fff00060fff2005bff8700a30079ffd10062ffb7fff3ff69ffee;
    mem[401] = 512'hffd0ffb7ffd300580031ff9e003bffccffe0006affa70069ff10ffd3ffdefff2ffe0ffc5ffd6008f002efff7005bff6ffffdff9a004bffd0fff5ff5fff84000f;
    mem[402] = 512'hffbfffa2ffda0034002bfffe003a0064003ffffc005dffa9ff62ff73ffb9006a0009ffec0042ff980058007b003affa0006e000d0046007b00b6009fff65ff7f;
    mem[403] = 512'hff7700810037ff44006affc7fff8fff0fff7ffe0ff85005cffa2ff4300aa0009ffea005c0014fffd0084009f00d000710058ffb20086004effbf0021ff9700e3;
    mem[404] = 512'h0015fff0fffeffc50011ffb7003cffbf0085ffe1ffef0038ff940002001a0087ff9affc60018007c0004008affd6ff6b00d7009cff42ffa6001b0098ff9800c8;
    mem[405] = 512'h0046fff8ff89ffab004c005b000cffae0073ffd70020ffc70082ff4800110068002effd5ff7fffda002e001f00d1fff9009f0000ffb3ff6fffeeff72ff650095;
    mem[406] = 512'h004100520028ff520087009b0012007dffee0026ffa1ffbc007bff61ffb70037fec900380026ff39ff96ffbe00770033fff10039ff7200da00380010004fffba;
    mem[407] = 512'h00b50048ff90ff6200570089006eff61ffdd0037007d00530144ffbe008600dbff7fffcc0070ffddffc10044ffca006d00b000aaffd9ff7dfff500afffc000ba;
    mem[408] = 512'h003cff8a005aff74ff74004dff4bff73ffa4ffdcffbcffefffa3005cfff20004ff7500960034000bffce005c005c008c0103ffec003c001e002f003b0018004c;
    mem[409] = 512'hfffbffb3ffcbffff000eff9e00770074ffd6fff5ffe2ffacffdfff80ffbf00e9ff92fff7005b000fffff0015fffd010d0019005c013c00090041ff580014000b;
    mem[410] = 512'h0039fff1ffd7fff3002fffebffd3ff69ffabff90ffec005a0016001700b60057ff8a005affe700550022ff99ff9efffe006fff690058001b001600850016002c;
    mem[411] = 512'hffa1008e005b00060016ffc7fefd0035ff8d00a0ffdc005f002d00650024ffb60013001dffaeffbd00420044ffbe0011ff8b0024ffa80022ffc20034ffe7ffb0;
    mem[412] = 512'h0076ff9eff81008b0001001100300077002affa40029ffe9ff650095ffec0073fff80011002cffcc0041fff4ffb5ffb200b1ff9600b40073ffc1006fff5b0021;
    mem[413] = 512'hffcdffe10040009bffe9ff68ffc90097ffa000390084ff430008ffaeffcdffb0fff7ffdfffa30098006affa500330023004ffff7fffafffafffcffcb00580066;
    mem[414] = 512'hff920022fff3003fff52ffe4ff9b006aff72ff920005ffb8ffd2ffa2ffa0ff5bffd9ff6f0073ffc00050ff6cffddff78ff96ffa4ffef004dff34007d00c6007d;
    mem[415] = 512'h000cffd90054ffcc00c9004200b80090004f0035ffb7008c0031fffdffc2ff5fff3cff78001e002c0086ff74ffd90071004effc6ffed00e1ff9d000f00f800b6;
    mem[416] = 512'h0003ff930026ffdb00d8fffb0082fff40011fff0ff3bff15ff5c002aff4a003cffe700a9001800d10092fff90029ffbcffdcffc1ffe0004b00690097ffa2000a;
    mem[417] = 512'hff61000b003bffe9ffad0056ff97ffdf00820054ffe1ff13ffb4ffc4ffbe0041ff92000fffcbffeaff9e0038006f0060000300b0003b000fffb1007600770038;
    mem[418] = 512'hff9c00070014ffd5ffd5004700270003ffc4ffaa00290083ffd90015001100fcffbe001500e5ffe90071ffa4feb6ff9affddffa0ffdfffceffdcfffa0015fffb;
    mem[419] = 512'hff8fffa90055002a000f00440031006a006aff890014ffe20000ffa8ff2eff5f0001ffefffe400500093ff9d0025ffddff30ffe90052ffe4ff9700ad001800ad;
    mem[420] = 512'hff4dfff5ff440010ffc0ffa7ffbffff8ffedff66ff6dff45006e0009006900140032ff76007dfff700adffc00050003c005a0014fff6ffdf0054ff9600160063;
    mem[421] = 512'hff6a007800510057ffdf007effcd00360080007c00910002fffdffbf007cffdaff5a0052006c0031ffca000ffff4ffc6ff95ff61ffde0064ffbb009a00a40057;
    mem[422] = 512'hff91002e003400160048001fffcd0014ff8100450010ffa70099ff7affadffcdfefa0076ffb8009eff87ff7dffa30032ffbcff9f00ba0064ffca0026ff58ff61;
    mem[423] = 512'h0055ffa8003b0088000affed005d003b0019ffdf0054ffffffb1006cff61ffa200b9ff7bffd700360035005afff300190028009b00bc004fff86ff7affcdff9c;
    mem[424] = 512'h000d00410004005dffcd004900260087003cffffff12ff820001003f009800baffe9fffc0022ffdb0027009dffecff94ffa70086ff86ff12001e0029ff60fff7;
    mem[425] = 512'h005e0001ff80ffd70042008bfff300410012ffe9fff4ffe2ffceff1f000a000c0009ffd50022009cffe9007affc6ff9aff54ffd40018ff260020ffd7ffb5003e;
    mem[426] = 512'hffb2ffdefff1004c001300310059ffcbff79008bff9c000eff39ffb1000700020015ff6f0053ffcf003effcaff77ffc6ffb40000fff3ffc8ffe8ffc2ff920000;
    mem[427] = 512'hffb5ff4bfff800a8ffaeffc6008bfff200880091002fff85ffaf002dffa0ffc7ff840029ff9f0072ff81006ffff3ffe1ffa100010041006effb1ff82ff55ffd9;
    mem[428] = 512'h007b002b001900aa0006fff2000e0017ff78ff3c00bfffacff1affc5ff98ff5bffa8ffc4002aff6600170048ffa4ff52008e0062008c0055ff43fffdff9d0052;
    mem[429] = 512'hffd10016ffab008e00480019ffd2ff1cff800061ffb70006ff24ff82fff5ffe400b1005300b40068ffe00089ff77ffbfffecff530023ff2e006bff87ffe0002c;
    mem[430] = 512'hff3cff9c001aff450043001f0032001300e6ff72ffe9001e0019ffbc0094ff3aff760065006cffe20049ffee00d1ffda002bff6cffc700200060007efe6f0049;
    mem[431] = 512'hffe9001fffc5ff830067ffc8ffeaff85005a0078ff7affd100220043ffd5ff5c0008fff9ff990022ffc60055ffe8ffcf0042ffb30014009cfff5ffd200220015;
    mem[432] = 512'hffa2ffd7ffff002400240024ff930012ffe30024001b003b00dbffbbffdeffc9ffd800ddffdcffb1ffb2001c0074008500ce00e80020003c001c001c004c0027;
    mem[433] = 512'h006fffaf001aff1dfffe00a3fe9dffa1ffcd0071ff89000bfff5ffc10086ffe7007300b2007dffdcffeeffd00061000d006ffffaffb3000b001efff7fffa002f;
    mem[434] = 512'h007efff5ff97fff700f400960018ffb00004009d0002000500630001ff8b001a00120020001b00420019ffe000010092003f0060ff4c0001ffba0088ffb7ffce;
    mem[435] = 512'h009c0092002dff8fffef0009ffe0ffa1006d0087ff71009b004d008800000005ff96ffec00d4ffb40051ffefffd200a3009f0021fff5ff67ff9bfff40044ff6a;
    mem[436] = 512'h0051ff6dff95ffba00820101004aff74ffffff71007100100020ffbfff79000400270007009bff1fffdf0057ffff00070005002800c90014ff9d00670004ffe2;
    mem[437] = 512'h008c0094fff7004effb1ff47001afff7ff560000000ffffeff58006100f8000500aeffebff5fffad002e0038ff7b008c00f6fff0012cff81004600850040001b;
    mem[438] = 512'h002f0025ffd40002002fff990049ff1a00e20069ff5800490004002c0041009300720062006bfedd002a008d005a001e008b0031005e006cffc8003f00900024;
    mem[439] = 512'h005cffeb0040000effbcff6ffff8ffcfff81ffc30059fff8ff2fffd5ffed0013ffc4fffafffeffa6000b000fffbc000a0077002e0070ffabfff80016ffc4ffaf;
    mem[440] = 512'hffb6ff42008bff840041001bffc1000e0009000d009fffcbffe5ffe5ff6affc9fff9009fffc1ffbfffcdffc400a70033ffc300310065000500a3ffe90017ffb3;
    mem[441] = 512'h003c003fff810037ffc100150088ff84fffaffc30070ff88ff9fffa5ff83ff93005bffa2ffb2ffe00014ff8200440021ffe8ff76ffde0098ffa9ff98ffe6ffc6;
    mem[442] = 512'h0002ffce001dff73ff65ff9cffdbffa7ffed00530037008cff40fff3ffe20023ffda00c2002d00330007ffd30026ffb5003a0058007bffd8ff77ff64ff95ffad;
    mem[443] = 512'hffb10028ff89007e00620051003500280099002d0066ffeeff5d001effd00042001c00060046000f001eff6efffdff3afff3ffbc012e00a30016ff950010005c;
    mem[444] = 512'hffc00089004f00480048004f00b900310082ff6effbbff96ffb9ffd5001800550035002400250061006b00c70064000afeb8001bffd4009c00a40027010900a1;
    mem[445] = 512'h0033002a0060ffbaffdf0015ffe1006d002aff82ff81ffd9fef4ffdc008a002d0018ffe400630057001cff5a00850002ffa10026ffa7003b00b0003f003bffe0;
    mem[446] = 512'h003affcbfffaffa4ffe900050056ffff003eff67ffb6ffd1ff7e003f002fff85ff43ff73ff86fff000b40007ff6a00000023005f0086004cff68ffb1001fff50;
    mem[447] = 512'h003a003aff46fffaffb20059fefdfffaff09ffc6ff9cff3e005c0014ffb80023003800b6fff8fff80018001300470066fffcfffc0067ffa8fff0ffe1ff8fff2e;
    mem[448] = 512'h0005002f002900a6006900570021005dfffc004bffd2006b00120061ffe2ffbb0006000700430025ff6cfffbffcefff5006aff82ff96ffee0008ff900005000a;
    mem[449] = 512'h004cffbaff620053ff950081ffc80069ffc7007e00250025ffe7ffb0fffe0013ffaf00e5001c0057fff70019000a0082ff89004cffb90091008aff7b0038ff73;
    mem[450] = 512'hffa2ffb0002f000a009cffe2ffeaffc5ffb300380007005f0019ff7e000dffa6001a0018005eff5effedffb300180079ffa30066001d009effc9ffa0001dffa5;
    mem[451] = 512'h007cffe4003bff03004d00e1fff1003dfff50097005cff87ff1d000affb8ffe9ffe8ffaaffbb0067ffa9000d0087ff9dff0affc3fffbff0e00b1ffb500bd0072;
    mem[452] = 512'h00b8ff5fffeaffe3fffe009fff9e0012ff66fff200b2003b0058fffd004f0039000fffe200120008ffaf0024003b004cff7cfff5ff98002a004bffdc00680017;
    mem[453] = 512'h0079ffcd006e002c002eff81ffe70056ffa6ffd7ff4d0046feedffab00830012002dff9a0044fffd005b0040ffb500a5fefaffa00055ffea0037005600f5ff74;
    mem[454] = 512'h00320048ffe100150061ff88ffd7ffde0047ff460094ffef000eff830089fff5ffb6ffb7ffea002d00650072fff20032001affbe00bafff0ffd600870019ffe8;
    mem[455] = 512'h0073ffba004a0085fff400ce0057ffa20095006f0097ff7aff51ffea0007ff83fedc005dffd4004aff8100aafffd00130043fff00043ffefffae000f003f0053;
    mem[456] = 512'h00b2000cffddfff5ffc800300063ff9dffea002000460071009dff6c00a8ffff003c003f0115005c00edffaa00500075005dfffe00a100a1ffba0011ff99009c;
    mem[457] = 512'h002d0039ff6dfff3ffc8ffbaffb7ffe4ffe8ff7eff75001a0067004c015fff9fffca000cffc6ffe6001effbfff72ff99000bffd7009b0036ffaa0059001e008b;
    mem[458] = 512'h0056ffde00a2ff920000ffaa00e4ff7a0043ff92ffff00b1ff65ffb30089ffdb0010ffe60070ffea00480020fff9ff7affd200930096ffd2ffa1ffdeff8d00aa;
    mem[459] = 512'hff77ffc7fff4ffca006e00d2ff89004a0048ffb000560085010700560090ffcfffdb00810060ffccffd5001d0011003e0056ffee00780032ff0d0032ffa400c2;
    mem[460] = 512'h002dff87ffc4ffc8007bff8c00b80057ff76ff67ff350001007cffebff85ffebfff0ff9a003fff25001000a0ffd00096005c0028ffebff67fefe0050ffdf0086;
    mem[461] = 512'h011cfff2ff86ffb3ff61ff9700a00009000bff7c006c00d7007dff5f002cffa5ffe10023ff8aff5ffff2000b00320014006800ea0082ff97ffc7ffdcffc20075;
    mem[462] = 512'h00faff8bffc70010000c0010ff70ff62ffddffc9ffda008dffb7ff8cffa3ff51fedcffec00710035ffb8007a0062000c00300030ff29001fffa8007e000a003c;
    mem[463] = 512'h0037ff3f00960048001aff530045ffd9ffe0ffc7ffd90002009aff0dff90ffcb000bff7a00e80037ff24ffa3ffe90006004500c10075ff3b009dfff7ff96ff92;
    mem[464] = 512'h00ffff96000bff28ffd0000bffc00020fffffff8ff93ff83ff9b001d00630064002800330018ff60009bffe90062015b0032000b003d004b0045ffcdffffffc5;
    mem[465] = 512'h00adffa900060042ff74ff81ff64001f0050005cffbc0033ffad005200750059fff0ff6500ca003bffe6003bffb8ffa5001fffa3ff9a004fff8b00320066ff61;
    mem[466] = 512'hffd700b3ffcb001afffcff7800a9ffbc003b009c00dafff6ffd7ffceffd20088ffe9ffc3ffc8fff5fffaffceffcb005affd9fffd006e0095ff8f0061000aff8c;
    mem[467] = 512'hffa5ffef002b00300009ff100002ff6c002600700058002cff6f00170047ffac0040ff7effc90029fed40000ffda00bf003600c4008bffe7ff83ffdefff30014;
    mem[468] = 512'hff7c0045ff27ffdcff97fffe0068ff8cffd400320035ffbfffd4006affe6005dffba0076ffa4ffe3004e0038006c004a0041003600380014ff4eff6f005bff53;
    mem[469] = 512'hff82ffd2ffb4007d0013000900330081006200820013ffa00026ffccffd2003e0021fff2ff9e007e001cff38003cffa9ff770037ffd9fff60028ff9f0087006d;
    mem[470] = 512'h0065ffcbfff900bb00c8ffdb00110060001800250001ffedffe4ff5dff5bff8d008fff7fff810035006f002b002bfff4ffbaff7900e5011c00160032ff950023;
    mem[471] = 512'hffcbffc40006ffedffbf00330027ffcfffe3ffae0026fed20001ff8f007efef9ff1d0025004affc5ff87ff3cff15ffc7ffabff51fffbfff000e0fff40063012e;
    mem[472] = 512'hff8cffffffd7ff95ffbefff4007a001c0056ffac0075001d00d7fffeffcb0001ffa4ffe8ffa80003008affddffdfffb8fff3ffc2ffb9ffc8ff8c000a001fffb0;
    mem[473] = 512'hffe0000affabffba00100045ffd100b0ff98ffdd0001ff8800000021ff45ffb90083001f0033ffd000a90049ffdbffa5003b002a006700ba001eff9b0042ffb0;
    mem[474] = 512'hffc8005100600003002e0018006dffc0fff6fffefff8ffdc0005ff31ffed0058006d001300770063fff0ffed002fffc5ffe7ffef0043ff43ffee0070ffaf0058;
    mem[475] = 512'hffb7ffbe005c0050ff83fff5ffc4ff96ff870075ffedff9400350081ff2e0012ff6c00cdffb80068ffdb004b001e008cffce0048003c0013001a0036008fffd5;
    mem[476] = 512'h00170052002e000f000d0053003000270071ffc400760015005fffdfffdd001cff8effd0007c001b008dffd4006f005900040049006a0009ffd2003fffc2ffb7;
    mem[477] = 512'hffe4fff90078fff400daffc3ffc5ff94ffc80032fff2ffc3ff6c0056ff890061ff0bfff70056ffd9ffd8fff0ffec00e1ffe7005afff9ffccff95006d0050ff8f;
    mem[478] = 512'h001500a0feccffadff4fffea00bf00bc0085ff90fff700a10027ffe6ff32001e003900750008007b005d00a200a7ffb100000067008d0058ffe10098002effab;
    mem[479] = 512'hff77fff80010ff91ff780084ff6fff76ffb3ffabffcf0007ffb80048003c009f00020035ff65fff5ff6cff68000fff0fff89ffb7ff4c003d0019ffeaff82ffbc;
    mem[480] = 512'h00c900a3fffc00070032ffcb00880007006e00550074ff62ffd8fed9ff98ffad002a00140046005400a5ffb80061ffb2007600560025ffb4ff9cff9e0031ffca;
    mem[481] = 512'hff920081ffd9001fff66fff2003500ed00a60079ffd4ffe4ffadffe2000eff82ff58005dffbb003900a1ff6effb4ffbbfffafff30037fff7004600a40077ffc1;
    mem[482] = 512'hffc5002a0071ffdfffaf0075ffcbffdb00c10056ffe5001f002affd400280074ffea0076ffe80005ff70ffe700220007ff41ff78000c0043fff2fece002fff83;
    mem[483] = 512'h0040ff1f0008005f009afff5ffebffc5008fffa5ff6cffbdff61ff1e007eff03005e001cfff5004c0079000200d0ffae0011ff08003dffa600cc007cffa200e5;
    mem[484] = 512'hffea0054ff42006a004cff980002ffb80053000f0029ffb200710050001cffb1ffd70006000f00e5ffe80071003d00af0037ffa50094fffdffacffee0001ffd4;
    mem[485] = 512'hff6fffee00250078008affc1fffbffa90006ff5cff68ffa600d9ff7e008affeb00740068ffe60082ffa3ff6600b9000fffeeff070053ff73008cfffcff3a003c;
    mem[486] = 512'h000f0069008800320052013cffd7ffaeff90ffb0fef60093005bffe9002dff94ffb200d300d7004400d8ffcdff26ff86ff8dff60ffe1ffacff5dffb10064001c;
    mem[487] = 512'h009dffeaffbd003900e7ffb800acfff0ffe20041ff110017004dffc400ac0033ff8c0040fff8ff99ffc0ffb8ffdafff7ffbdffd000d7006800b90180fff10072;
    mem[488] = 512'h006d0072002b000f002c001bffbdff45ffc1ff97008affd500970040fff7ffc90062ffec0019ff630015ffff0110ffc0ff5b006fffe700c70070002d0006009a;
    mem[489] = 512'h00c2ff5c0049ffadff6f0039ff65ffd0004dffd3001800660043ffa6fffaffc50043ff360050ffde0002009700d100640060ff650041004a0010008800050052;
    mem[490] = 512'h00940086ff89ffc2ffe1ffd600ecffee003e0048ff38007f0086ff7bffbcffc00062004effe7ff95008000110028004500070029fff2003effa4ffcaffccffe5;
    mem[491] = 512'h00cc0049005b003affb7009cfff7ff48000bff95ffd7009cff74004f00460004003f00120051ffe3ff5801180047006a003c001000a4ffee0048fffe00b8ffb4;
    mem[492] = 512'h000c0053ffe70006ffbcffba000b003b007bffbc00280000ff12000bffdd006dff610030009d004dffbdffbb0061ffc3007ffff10034ffa9002eff76fff1002b;
    mem[493] = 512'hfffa0009ffb2001f0058003e0007fff7ff9dffa0002400150015ffe100d6ff45004e00490009ffcc0037ffaf0023ffde001cfff200220034004eff56fff8000c;
    mem[494] = 512'hffa20059002dffc90074ffc000aa0017ffbeffd90042ffd5000effff002500170010006effffffe8002b003afff0ffb60049ffd2009dffb3ff80ffb2ffaeffc2;
    mem[495] = 512'hff75ffce0055ffa6004dffd0ff16ffa00024004cffbfffc8ffddffe000170034ff5600cc009effe801070021ff620052ffb8ffef00b8001ffffaffc0001ffff7;
    mem[496] = 512'hffe5ffccff9d00df007a00370067ff83ff7a000dffe7ffd4ffa20035ffdafff7ff940006fedf00f3000fff820087005e0095fffe00110094ffd7ffa5ff7affd8;
    mem[497] = 512'h002c000dffa70001fffe0021002f005eff9eff63ff9bff1b0018005d0064ffee001800b7002b0016ff86ffcf00510030fffeffeb00510051ffcdfff6fef0ff95;
    mem[498] = 512'h004a002c00100039009b000100daffe90010ff49ffaafff5ffb900510000ffe2ff51000fff8b000800460066ffe0ffadff6e000bffcafffdffe900230024ffa4;
    mem[499] = 512'h0080ffcbffdeffd30001002c008affeeffd8000800d5ff46fffeff85ffcfffc400b9003a00030032ff8100df003b003fffdf001dffa7ff42fffffff6ffef0021;
    mem[500] = 512'hfff9ff4d008affc30052ffb3ffe9003fffa20018000f0088ffdb0039ffbc0012ff6b00430004fff60019ffb4ffcf000d0059ffecff750008ffb70049ffef0039;
    mem[501] = 512'hff7effee00770019fff0003aff750060ffe200650023004eff62001e00490039000bffa0ffffff67ff91ffb80051001f00000020005affaeffc4ffad002cffbe;
    mem[502] = 512'h00360083fff1ffefffe00012006f0010ffbf001e007dff78ff77fffc001000380021ff28ffd1ff35003500d7fff50012ffe9ff7c0002001dffdeff6effadff50;
    mem[503] = 512'hffbf000900b1ffe7ffcb00090085008300690089ffa0ff7affbaffed0009ff200021ff6dff8effec00080058ffa4001f0107002b0105006d00270068ffb4ff80;
    mem[504] = 512'h0100ff3800370105ff7900230015ff8e00130055ffdcff90fff3ffd500f8009f006800170040ffe1ffd900c2ffe4007dff9bff8d00100014ffe2ffa7ff690144;
    mem[505] = 512'hffcb0007004f004e0004fff1ffbf004f0021ffee002200210075002c0053ffd5001fffd900b7ffcdfffc0037003b00160030ffe000030028ffe5000c00330026;
    mem[506] = 512'hffc9001e0009fff0ff76ff97ffb20085ffaf005d0056ffa9ffca001a00750001003c00a1003d004700340074fff7ffcc001c00350005ffe5ffe8ff8bffa90074;
    mem[507] = 512'hfffeffdc004600660043ffb1004c00ebfff8ffaaffe6ffd9fff00084008b00c5ffb50058ffb9ff74ffc8ff49002200780031ff8affdc0076ffbbffe4ff2b00d9;
    mem[508] = 512'hff85ffb8fffbff7d0052ff40002cffa8ffc50000ffcfff8affc5ff89002500a20026003eff37ffe8ff94ff82ff98ffe4008cffa30006ffe8ffba004fffc10032;
    mem[509] = 512'h00030052fff0ffb6ff62ff540063004b00a2ffd3ff32ff56ff950049ff92fff7007c0015ff3f0002ffedffbfffb0002fff7c0044ffd8003effd6001dff99ffeb;
    mem[510] = 512'hffb6006cff34fffc00450045001a00940082fffb004d0012fffb0055ff370006ff9bfff5001a0040003e008b0039ffb1ff58ffa3003f005c004dff7e00960014;
    mem[511] = 512'h0071000200160032000bff99000b003eff440002ffb2ffe4ffc50017ff9000050064ffb1001800e300ac009800150013001f000dfff60003005bff8d000700ee;
    mem[512] = 512'hffceffa300520082fef6fff3fff4ffd200c50077005e00150074ff810026ffc5fff1ffcd006fffec011300340049ff50ffcf001affbbfff30044ffd9ffe6ffe3;
    mem[513] = 512'hffe8ff6d00430032005e006b0064ff62ff7aff2c0004ffe1fef900ab00c6ff6a0040ffcaff73ffbbffd10083ffb10047ff210005ff67ffaefff70045ffef0050;
    mem[514] = 512'h0057ffbb0053ffd000eb0022ffb2003a004dffe2ffafff81005cffc1ffe9ff25ff8cfffc0039ffdd0042ff29008e0047ff8d0026005cff77ffc4ffc3ffb9004c;
    mem[515] = 512'h005dffffffd9ffd7005a001bffa0000c00390021000400540032ff07ffa20065002e0022009100a2008eff91000effcbffb9ffb1006d001400d4013eff93004b;
    mem[516] = 512'h0022ffffff87ffe9005fff400022ffb300dcff6cff71ff9b0045fec0ffe1ffba001d00a3006bfff0008c00330040009dff730078007eff8500160008ffc50047;
    mem[517] = 512'h00d7000c0021003dfff800d10053001afff4ffb0ff64007f0033ffbdff3f0058ffd1000700f5ff97ff11ffe6001dffdfff63ffdb003b0075001cffb90064ffbb;
    mem[518] = 512'h00d200040038ffbaffb300bf0092ffecffd8ff42ff730073005fffef003dffe50097000ffefdff78ffa60008000cfff7006b00f7000200d2ffd7002fff8affc9;
    mem[519] = 512'h006bffa3ffa6ff52ffed001fffee001a0018001f003c00280012ff7c0070ffcb006aff7200580027feceffa10018010affcd002d00c5ff79fffaffab0045ff1e;
    mem[520] = 512'h00840008ffd2002dffd9000b0037006b003f005500190037ff530018ffd6ffbfff76007affe8ff8a00730019006a00140009ffe3004f00260051ffeeff9b0061;
    mem[521] = 512'hff78000cffc40039ffeeff8e00480077fffa0052009cff330021ffa6ff5bfff70042ffb200370004ff76ffd2000afff20046000e00a9ffc70005ff5cffebffc5;
    mem[522] = 512'hfff700dd003afff2fff200a10046ffd6fff80052fff3ff900020002b00440053007c00be000400000018ffc50055ffb9001affdd006effd2fff500a50017ff70;
    mem[523] = 512'h00810026fff50055ffee00a0006a00a70000008efff1ffaeffec00a0ff6affd0ffd5ffc7ffa1004d001bff5b0088ff6cffccffd8ffe4000bffb20079ff960019;
    mem[524] = 512'h0040ff53ff9cffac004200860037ff97ff55008bfffbffac001b0030ffd3003bff87ff94fffbffd00011ffae0021ffd8001bfffb002c00b9ff8d000effc60057;
    mem[525] = 512'hff60ffd20068003e0073ffbdffdb006d008d001d00c1ff44ff940062ff8bffadffdb003200a6ffb9ffd7ffd5ffcd001effeaffe9fff7004c0042ffe0ffddffcb;
    mem[526] = 512'hffac009d000aff67ffe5ffbb00ce001dfff200ceff5dffefffdf0021ffaf0074ffd2003d00860090008a001affd500d2ffe2ffa6ffea00d2001fffd8008cfff8;
    mem[527] = 512'h00a500670015006a0096000d009d0123ff7b0027ffc1ff9100140020fffcff58ffd6001dffeb000effbdffa900140065006e00a30050ff9effc7000f0034ff99;
    mem[528] = 512'h005affd0003c000c0052ffc1ffd20059fff60014ff8c00230022ff58002bffa7000a0033ffe4005b0068ffe5ffb3ffc70048ffb10047ffeeffe8ffd4006f000d;
    mem[529] = 512'h00400032004f0029005afff200c30081ffbf0021ffc90069ffafffe9ff730044fff3ff84003b0013ffb3ff9a0026fffe007bffac000f000bfffdff95ffd30034;
    mem[530] = 512'h0069ffd0ff160008ffbc001affcdffd5004000440014004a0067ffcd001e0026ffbaff76ff36ffd6002bffffffa0ffcdff6effe0ff8bffc00002000300770015;
    mem[531] = 512'hffb9ffdd006dffcc0032003800920030001400b4ffbc001aff62ff9b00840012ff5dffbbffd7ff36ffa0ffcfff9c00830044004dfffdffd5ff8afff800800063;
    mem[532] = 512'hff9c002dfffc002200440048ffe8000400460020006bffe6005b001c0046000a0068000600c5ff8dfffb0076ffcfffb0004dffbbff7b007f00350024001c008d;
    mem[533] = 512'hffa7ffa90065005b001e004dff9400a00027ff85002500160002ffce0022002900580019003bffcbffc7ffac008c0016ffbd0003ff9b001e0033ffc1ffa5000c;
    mem[534] = 512'h011a006e0027ffae0025fff1001f003100920006003fffb2000dff3e006d002a001cff80ff7400070034fff30077ff810041ffe3ffcfff320069008400290037;
    mem[535] = 512'h00410038ffd10035ff9f0072ff76ffa9009900570008ffbdffbc007c0047fef7009800fc0041ffb9002d00d2ff9600630047ffb9ffe1ff8500640002ffbeffca;
    mem[536] = 512'h0018fff90052ffd0ff8dff650036002affaf0000fff5ffb9ffedff81004800a10062ffc5ffd9ff9effaa004eff77003800540042001dffa8ffdfff7f0079fffd;
    mem[537] = 512'hfff4ffc4ff87ff6bff840018fff30020ffd10025002a002a00a90030003c0015ffdc008d00640037ffaf0011000e003f0099ff340006ffd30066fefbfff900b0;
    mem[538] = 512'hff05001bffa3ff82ff32ffba0030008e00a4ffaaffa0ffbeff6fff4f0072000000610015ff6efff1ffb300ab005000a7fff6fff20030006f000ffeacff9fffdc;
    mem[539] = 512'h0066ff73001afeebffd2ff48ff520089ff950085fff7ffa40063ffedff27002d0021003100a7001e0038ffc20012ff54ff8700270027003300d2ff76ffd60031;
    mem[540] = 512'hff48ff460024ffeb000d001e000fffde000a0029ffaeffde00600019fff2ff4affe2001effe800e00035007f007dffaffee500460015ffcb0023ffc0fffb0097;
    mem[541] = 512'hffcbffbbffe8ff94008cff5dff3700e5fffeffd7ff92ffc200620026ffd8fef0ffc40023ffc1ff87ff79ff99ffb5ffb2fff5ffbe007c006b002e0027000600b7;
    mem[542] = 512'h0054003effb000a2005fffc0007200b2ffeffec7000dffd4ff95000500020061ffbeffa300b80073ffb4ffe1005fff81ff4d0052000cffc6002e0031fffb0097;
    mem[543] = 512'hffa6005f0059ffc3008f004effbd001a006cff5100900072ffe5fffd00310002007effcfffbbfff1ffcaffe50005ffbeff2e00520025ff9b00b8006d0023005d;
    mem[544] = 512'h002e0025ffde00590045003b0051002a0017ffbfff3b009e00160057ffb0fff3ff34013000620053006f00e700f1ff9cff9f0011000f003bff3dff9fff65ff94;
    mem[545] = 512'h0043ff75ffaa0020003cffc4ff42ff7200110039ffae0056000cffe6002a0021fffaff45007affff000e004cfff3ff92ffe3001b0020ffa6ffa50024ffea0059;
    mem[546] = 512'hff4a0071ffc8ffc301210041ffbd0024001b008eff78ffcbffedffdaff9dff93ffad007f003cffacffe10023ffcf0017ff52fee8008a0060ff42ff610059ffc8;
    mem[547] = 512'hff6c002f0019ff9000060086004affdf0073ffc90023fffd00240006ff770021ffae0056ffe2ff32ffb30007fff7ff8e0058ffa1004300010029002fff880054;
    mem[548] = 512'h001b00120005ffa6fff8000effebffd2002d0098ffa1ff460104ffc100000084ff8100590033fff5ffa4ff83005b000cfffe000200ad0085ffaffff1005c0083;
    mem[549] = 512'hff6bffaaff67006a007b000300600029ff780006ff9bfef00002ffe1ff5c0118ff68ffe2ffc2fff9ffce0054003e0007004d008f008c001effdcff6a0071ffb4;
    mem[550] = 512'hffb3ffbe004cffdb0092ffe5ff4700faffa9ff880090ff7fffe1ffc300040069ff3b00130054ff42004500150050ffb00011ff8e0026ffec005e0058ffd600cc;
    mem[551] = 512'hff8800170028003a0005ff6fffd70058002400d100670067001e0051ff8d00c4ffea005dfff4ff77001affe300d7ffaf000cff76feecffb2ffb1003cff660010;
    mem[552] = 512'h0013ff97ffdd00f3ffd8ff2900200024003000d30088ff92ffcc00810061ffff01000050fff6ffa30046ffae00330078002e0011fff5ffd50003ff81ffcb00a5;
    mem[553] = 512'h00080081ffd6ff33002a002e0004009affc0ff07002f001dffa10010009200b7ffd70010ffeaffe0ffe4ffa7008dff8c0061002d0052ff6cff9bff7affec0000;
    mem[554] = 512'h003fffe600eb002affe8ffa2008e00210031ffbfffe6ffa00095ff2cffea0021ff29ffe6009c000eff970044fff2ffe200dd0075fff3ffd90020ffee00000017;
    mem[555] = 512'hffc1fff7ffeb004b000affe1ffc90060ffd60080ffbaffc70029ffddffe3ffc4000e0011ffb6ffe8ffc40013ffbe001b00230075ffeb0005ff37ffcaffb1ffec;
    mem[556] = 512'hff6d00630012004e000e00790070fff2005500d000420084ffc30020002bffceffc5005dff83ff45001fff81ffe10070003f000c0018ffffffecffa7ff66002e;
    mem[557] = 512'hffe0ffa10001ffbe0026ffeaffc9000e003a003e000a0081000c009bffd7005cffe5ffbfffd2ff560031001b0046ff8d0006ffa9ff8fffed0060ffe00045ff28;
    mem[558] = 512'hff8b0005ff9000990079ff950049ffdc004fff9b00e2ffda00a1005eff3100320019fffb00b6ffd3ffb6ffeafff30029009700240033ffe70036005fff990047;
    mem[559] = 512'hff98ffefff220049004f0004fff2ffb7ff3b000c003c005fffdf003b004f005aff550060ff84ffed00cfffe5002bffe4002e00ab005a004f0035007affdaff75;
    mem[560] = 512'h00490057fffa001a0024ffda003bffc4004affe2ffe4ffc4ffd2ff8cfff800040001ff6600320051ff0cffb5003d0081001e000a00180035fff8ffedfffa0031;
    mem[561] = 512'h00710005ff560041ff2d005fffba00b3003aff3dfff10004ffb60057ffe20094ff68ffc50064ffea0023003bffccff8fff99ff1fffedffd3ffcf008a007c0076;
    mem[562] = 512'h004bff760065002b00e3008b0038ffb4ffedffd5ff3a00d4ffe6ff67ffe8004dffdf0083ffe6ffe5ffc3ffe40027ff660040ffedff63006e0063007f0026fff3;
    mem[563] = 512'hff8d001f004effb5ff6d00afffdc0003fff5ffbb0094004b002b00370012ffad008eff750022ffe20055ffe800a3002a0050ffd4ffe000660014ffbb00840073;
    mem[564] = 512'h0081002000aaffc3ff8f000eff1e00510068ff9eff820054ffff0079ff56004effa4001cffd900720031003effcd0009ff83000dffcf004e005affe40049ffb1;
    mem[565] = 512'hffd2ffe4003cffffff93ffb100270030ffdd0020ffb00028ffceffe7ffb8ff98001f000d0059ffba00a4005000330042ffcdffa800000011006c0061ff920083;
    mem[566] = 512'hffb5ffe3000e001c0068000f004e000fffbbffde0049fee8009300f70013ff2b0016ffc2fff700080018ff8bff7dffd30005ffacff2cffd6ff5fff3dfffa0024;
    mem[567] = 512'hffd10035fff10004ffbcffa8fffe0029ffe8ffe40075ff1a00910036ffa2fff7ff80001000350073000400340066ffab0046ffceffb6ff67fff3fff700320041;
    mem[568] = 512'hffebffef012d0066ffe2fff4000f006f0091fff9fff3002d005e00770001000000ceffb2ffe60011006bffa90021ffe0001e0024fefaffa9ffb8ffdf0074003d;
    mem[569] = 512'hfffa0019ff90ffa000400059009600960039002e00000038ffd7ffebffd6ff230008019fff8f004dff98001bffffffe8fff0ffb0ff780022002c0029ff94fff9;
    mem[570] = 512'h00150049007f002400380006ffbf0069ff980078004b001b002000400013ff34ffa1ff7500220049ff69ff940029ffbdffd300190021007effd10022009a004d;
    mem[571] = 512'h0068000600720048008b0038006c003b004affc2ffeafff3008effd8ffbaff6900b8ffcd0034ff90fff0000d00300033ff67ffc3001dff8cff77001fffeb0066;
    mem[572] = 512'hfff800bbff1d0068fffafec9ff27003f000dff76000c008dffd7fff5ffa7ff9e00b5ffad00a900160035ffe40169ff88ff85006e0092ffd40096008a00aaffe5;
    mem[573] = 512'hffe40026ff84ff990002002a001affca00a5ffd40031005a0095000bffec0003fff00063ff87ffe70092ffebfff10018000000590040ff8a009bffdc0058fff3;
    mem[574] = 512'h00690089fffeffe20065007fffbaff77ffb4fff100590006ffb6ffe9000300390097fff1002c005cffadff3500c6003d0072ffb0009b005dffe4ffa3006f005c;
    mem[575] = 512'hffa40003003c008500c7ffe5ff3bffaf0006009fffa60037ffd3ffe1ffbafff9ffec000e0070ffe50023fff900450053ff79ff89ff51000cffd0ff8d00a5006d;
    mem[576] = 512'h006c0011ffb7003f009f004affaa00570059007c0028fff2ff4bffffff9c0026ffccff730013ffbd006300160007ffb6fff6004b005affcaffbdfff0004cffee;
    mem[577] = 512'h0004001d0001ffcc0059ffffffa0fffdffe3001fffc8ffd00019002400300059ffe4ff8cfffe005b0041ffc600a1ff70fffbffe50067004fffdbff8affefff99;
    mem[578] = 512'h006400250035ffd400d9ffa2009dfffbff5a00ba004f001c00490023ffd1ffcb001100290072fff6ffc1002d0056ff3bffd8ff27ffd5ffe70065ffc7ffac0049;
    mem[579] = 512'h0015fff30033ffdeff760028ff3bffddff9effdaff9fffa1ff82ff9400520021fff1ffb60061000800140043000afff400030009fff7fff2ff2b002f00590040;
    mem[580] = 512'h001effa800560060009d000eff860074000e0113004f001d0023fff6ffa00027005f003d008aff86ffc4001d0023ffbbffb0fffcffa1ffd60042ff75ffaf0079;
    mem[581] = 512'h00af00c20008ff890042ff9affb70083ff9d0005ffa0ffad00450004ff84ffc0ffc9000c00a70049ffe60017004d001f001c005fff74ff5f0029ff9f0063003a;
    mem[582] = 512'h00020005ffc60002ffb8ff63ffc50015ffe9000effae001bffec00f9003fffe2ffe9fff0006a0046003bffc8ffd7ffa60034ffcfffceffe2ffc8003600d2002d;
    mem[583] = 512'h001c00be001e00a3007f00110101fff5ff9afff80004ff1d0048ff780053ffbb00090073ff90fff2ffe60003002aff7d005fffbeffe700180016003eff87000b;
    mem[584] = 512'hffa100d2ffcbffd5ff360026001f0015ffcf00050015fff70031ffa2ffccffcffffa00880031004d0098008a004cfffb001f00d5ffa9ff80ffe9ff4300d4ffcb;
    mem[585] = 512'h0056ffa5ff890091ffa10092000affc4ffcafec7ff8eff6affad003cff94ffe6ffb4ffbd0018ffc3ffe7fffeffed00af0054ffe2ffb5ff82fff100bf004cffd0;
    mem[586] = 512'hff92ffd4ffc0ffddffa4ffee0045ffc5005200220006001afff2ff75ff9cffc8ff66003efeec0043ff91ff7a000effa50005ff50feedffceffbeffe5ff910003;
    mem[587] = 512'h005000c8007dff94ffacffa5001e00380005ffd30062ffa4000efff9ffab000000570045ffc9000d0031ffe4ff91004fffa8ffabff8c0047ffeeffe400930019;
    mem[588] = 512'hff7cffca0086000afff200080085ffdd000c00aeffcbffc4ffa5ff88ffb90082000cffa4ff8affea00c3ffa0ff96ffb9fff9009f002d002dffb5ffa300590076;
    mem[589] = 512'hffe4003eff750036ffc60018ffc200ab00910002ffc2002efffc009e005d004b001700e6005cffffffe20019ffd9001b0009001f01540061003bffe1008e00d6;
    mem[590] = 512'hff7aff9c00b1000affccffe9ffe1fff9ff500084ff9c00360090ff87ffce0036ffebffe3ff3f00f0ff97001dff7f00c9001e006eff960076ffe6ff85ffdf0058;
    mem[591] = 512'h000cffd300430050fff1ffc6ff65001c00b0ffc50036ff97fff80016002d0047ffe40068ff8cff770014004e00320053001eff5b0091ff7aff4b00240076ffa8;
    mem[592] = 512'hffd00020ff90fffeff32ff30ff620003009200220065ffb9001cffbc0011ff90ffb7ffebffc300290010ffcc0015ffdcffedffdfffb1ffb00009ff830042007c;
    mem[593] = 512'h0079ffd80022002bffa0ffe60019ffafff0cffd4fffe0026ff620020ffec0033ff9b0057ff9dff72ff3affc10002fff0ffef0022ff32ff76ffd3ff8200d5ffce;
    mem[594] = 512'h00770040ff86ffbcff89000f0011006c0044ff9a005a00b5fffcfff0ffd7ffa4fff20015ffbc0042000900040090ff45004f0034ff8bfff9ffb100cf0066010f;
    mem[595] = 512'h0027ffa20022000eff820020fffeffcb0102005e003c004c0079ffd2001bffc9ff7a0031ffe0002dff3000b90020ffdf003700430031007b009dffddffdbffef;
    mem[596] = 512'h00080003ff1b003000330048ff7e006d002afff20030ff8b00ddff6c0035006b0016ffe6fffd00570096ffc80011ffa8000b001fff75006effd4ff5800420092;
    mem[597] = 512'hfff000abff81ffe8ffaaffc8ff620021ffbfffa3ffb2ffddffa2001cffb50040ffec00160052003cffd2000f0035ffc500890083ff80ff8effce0083ff5ffff9;
    mem[598] = 512'h005e0088ff30004fffdb006affefff72007cffcd0074004affbd00780032ffd9ff7e009d0105001f0021001d00780028ff2c0029002100b00113ffddffde002f;
    mem[599] = 512'h000100780040ffdc00580051ffbc007f007d00c7ffee0033ff4a008bff83fed8ff730076000f006f003e00060053ffd9ff68ffd9ffdcffa400c7ffc00022ffea;
    mem[600] = 512'hff4c002e007cffd80131ffccff40ffddffef0084ffebfff400350021ffb3ff9affc3ff5a0058ffec004b001a0056ffcdffabff5affd6ffa6006c00730083fff9;
    mem[601] = 512'hffd1ff9bffd6ff97013c0041ffdc008100330011010cffd300500028ffb7ff7dff64008a001e0007ffcb00bd0010ff72ff57ffb2000a008eff960029ffadffe2;
    mem[602] = 512'hff6400c1ffb7fff0005d009dff9f003b007f004bfee0fff9004100bcff21ffa600170024000cffb6ffbf005bff9e00d100c5fff9007100200056ffda0055002f;
    mem[603] = 512'hffe90074ffda000400440049ff64000eff91ffebffceffbdffb6ffe8ff5b00cc001a0016fffe011dff7effc3006fff47ffcfffe60005ffb4fff5006b00180011;
    mem[604] = 512'hfff0ffd1ff8affd80057ff84ffea009ffffaffed0080ff0affb0fffffffd0057005d0041ff4c00240033fff4ff5bffa3009500640068ff8dffcfffd7ff8dffeb;
    mem[605] = 512'h00b60036ffb9ff85ffa20048ffbeffccff33007c0044fee9ffccfffd007600cb006c008fff99005effa7ffdb0061ffe600970019007400430033ff4cff68ffcf;
    mem[606] = 512'hffd200500001002f000a004dfef50027ffc700060005ffde00a2fffd0003ff88002affe2ff9dffed0019006300b3ffac011000070039ff2aff47ff8effa1ffc0;
    mem[607] = 512'h0010ff5f002c001c0033ff54ff2e00a7004100130095ffdc0016ff58fff1ffecffefff9affd30008ffdaff72009d0067004effeafff50046ffaa003cff9700c7;
    mem[608] = 512'h0079004bffae00690055ff5900700062ff94002fff4efff90094ffa000810029ff9cff99ffc1002aff5b00c9001cfffdffba001a002efff200240048ffe9fff1;
    mem[609] = 512'hffa8ffae00b5ffa70052000d006000daffe400a9ffcb002eff80ff51fffc00540036006aff2f0038ff94001e0049ffc8ffc8ffb2ffcbff9fffd9ffc9feefffcf;
    mem[610] = 512'hff7c0064ffb900a70028009f002a0084ff4bffcc000b007100fcffe8ffcdff7effb6001900790049ffb200ab0047fff5004ffffcff32ffe0005600a4fff1ffd7;
    mem[611] = 512'h003eff870015ff9fff990001ffa7ffd1001fffcaff96001f011b0000003eff60007000420044ff78ffbdffc90016ffc8ffe0ffe000f6001c00e00005001cff7c;
    mem[612] = 512'h0009ff9dff2effb100cbffd7001d006dffdc004000230055ff780084ffc3000eff820067005cffd7ffd700caffe6002b00370081006fffcf00640033ff5f003a;
    mem[613] = 512'h0038ffb90005006a0065ffd8ffcf000cfff500870066003fffd9ff8700b5ffc3fff8ffcbffdf0071ff2ffff5ffdd00700074fff8ff35fff0ff40ff2c00010003;
    mem[614] = 512'hffceffa7ff99ffe8fff3ffb6ff58005700d6003900a60029ffaa008fffd4ffe400f20012004dffd40012004d003dff9b0004ffe30025ffc30016ffa4ffa000ad;
    mem[615] = 512'hffe300320045fff7ff920016ffaeffcf00820036003effd7ff96fff8ffb9004affe0ffc5ffab002dfff2ffb8ffca0032ffbaffcc0074ffea003fffc5006e00e4;
    mem[616] = 512'hfff4008f001a003ffff4ff90ffa3001dffb7004f0029ffeeffa60087fff4ff3a00ae003d0004ffbdff8900080077ffc4ffdc00100058002900e6fffd00a40000;
    mem[617] = 512'hfff700d7005bff8200c1fff9ffb8ffa40047002a0015ff9b00010043001a002a0074fff3ffde007a0016ff53ffaa004b0047ff950020ff68fff2ff8bff93ff62;
    mem[618] = 512'h0025ffeaffd700420037009effe200390004ff77005500860012fffb002affdffff1ff570023ffa0ffe3000a0041002700de0018004bff8cffd1ffb10044ffd8;
    mem[619] = 512'h0011004d003effa3ffbd00020042ffb0ffeb00ab002a00430020ffe4001c0012008eff290010ffbbff78fffbfff30025006f0035ffc7ffcbff9c00740033fffa;
    mem[620] = 512'hffc3ffd5ffbb0043ff72ffe3ffb500190087ffd90037002aff100021ffd6ff76002c005a000bff7a0077003bff80ff82fff800610015002b002d0091ff8f005c;
    mem[621] = 512'hffc0fff10023ff6affb70003ffff0038009100300039004d00100098ff3900aeff69ff6c004fffac002dffb9000d002200d4009100bdff2dff63ffbb007eff36;
    mem[622] = 512'h008effefff9fffb800c40093ffe700b9ff76ff840083006c00070035002fffbf0070008effcd0021ffc2ff79ff530015ffe90011ffdbffbf000eff7700960052;
    mem[623] = 512'h0105009cffb200a5ff96002e004d00ad004900a300070067ffff0039ffd6002a005afff50035006fff8aff860026fff3ff83ffecff80003bfff0000a00790008;
    mem[624] = 512'h003a0039ffdeff44ff8d00b9ffff0077ff560031ffd6ffeaff4f00280005ffd6ff76002dff4a00540001000100260029ffbf00730083ffdf0089ffef0014005c;
    mem[625] = 512'h0060003300280083fff3ff07fff800a3fff80066004bffc100aeff98ffbd008e001dff3dffe900670043ffe8007dff6e004b003b0013ffbb0038fed5000700ab;
    mem[626] = 512'hffd6ffadffafffdcff91007e007500b900700040006e002c0000ffc100790024002a002b00d6fff0ffd1ff90ff75ff720007fffbffeb00c1000bffbd00b10029;
    mem[627] = 512'h00ae00740005009bffe9ffc9ffc600a8ff0bff4a0002ffcafffb0001ffe7004fff70ffa7002300da0037ff6200fa0070000dfff4ffe0008300d5008e0007ffc0;
    mem[628] = 512'hff3bffa5ffc00032ffa6006dff6400b2ff56ff82005b00690081010e0074ffc50069ffd0ffd4ff54003d002800bbfff50062006f000000240043006600b3000e;
    mem[629] = 512'hffd8007cff9efffdff7200490035003bffd2ffb4ffd6fffe0011ffeeff84002a005a0005004bffe60094ff4a002affd50051fffc00d8ffd7001c007cffe7002e;
    mem[630] = 512'h0009ffb1ffa9001cff89006dff99007f0059ffbeffaaffc400630066005c0039ff910041009cfff8ff78ff64ffe8ff86ff9500ad000aff87fff6000a0019ff93;
    mem[631] = 512'hffd0005d001cffdeffd8000a0016ffac0035ffe20059ffbdffd1ffb10041007afffdfffc00930032003f001d006c003e007700620029001f0075ffe2ff83004a;
    mem[632] = 512'hfffa0042008cffe200260022ffa8ffe5ffdeff84000e005d0077ffd70035ff9bfff9ffc6ff38003dffd3ffc300cdffb5ffeb00affff1ffca0095ffd3ff920000;
    mem[633] = 512'h00480094ffb00016005f001cffbb0064ff64009affebff07fffb00d9001dff50005d00310050005affbdffee00590012003e0072ffccff5dfffcffa700550005;
    mem[634] = 512'h003f00250023ffc7ffdbff5aff2e002a00640085ffe0ff62ffa0fff70007001bffe40082ff79ff8800a60098ffee005400150005ff8f001b005affa9ffd5ff78;
    mem[635] = 512'h006dff48004a0061005efffeffb5ffd0ff6bffa50015ffc9ffe5ffd0ffb1ffbfffa6ffdcff89005f0018ffea0003fffe00a70044ffdcffa400bbffb300730078;
    mem[636] = 512'h006401150047002affcaffbb0078003f002300aaff72ffcfffe7ffdc0005ffe00004001bffce0009ff83ffd8002aff94ffc000b4ff7b0063ff96ff2ffff6002b;
    mem[637] = 512'h000affb0ff810028ffbb000d004affa8fffdfffeff5fff51ffd6000dfff3ffad0049ffbdff04ff8b000dffd00048006dffde0044007f0046ff5d000aff77ffec;
    mem[638] = 512'hff41ff6600a2ffbf0001ffa2fff200440076003afffc001aff650010004cfff300f7015affe7ffd5006dffb9002bffa5fff5009dffe4ffc9ffebff92000d003b;
    mem[639] = 512'h0003fed200880015ffe70079ffcf0005001bff57ff37ffb1010b005effc70081ffbdfff600200024003100ba00a20026ffbeffe6ffc90000006fff75ffc4ffd6;
    mem[640] = 512'hffe7ffb3ffbe002200590055fffefff6006e000b009c001fff84001d00430069ffe2ff160074fffa0034006d004effe70018ffe30002ffa9004e00c200380077;
    mem[641] = 512'hfff0ffbeffedff7cff60fef6001effe8ffe2001d0027ffae00340081000cffad00c5ffeb0037ff97ffd50015ff5cff7200370071ffa5fff9002f000c00490074;
    mem[642] = 512'hffa0003e007a0083002dffe90041ffe20063ffa10026ff9a00abfff6002eff95ff8b00caffeb00e1ffe3ffcc008bff23003cffbfffda003a0015fff900e6ffda;
    mem[643] = 512'h00a8ffd8fff90043004fffebff9cff240062011d00240016004900090021ffd1ffd6ffeeff68ff0d0011ffdfff92ff670041006a0088fffb000500d6ffdb0080;
    mem[644] = 512'h0039006c000e0085ffd0004affef00820009003b008700a9ff210047ffe6ffb8ffa0ffddff88ff7fffc3000cffd8ffc7002fff0aff7eff3dffdf00c6ffbdff75;
    mem[645] = 512'h0066000e0084ff4b0076006ffff0ff9effeeffc80051ffbb0024000e005f004b00ec0016ff5dffc4ffce0029ff6c006bff5d006cffb4ffe8006d00930004000b;
    mem[646] = 512'hffecff97ff59003000c1001bffb3ff71ffc200400082ffe70044ffdc0095ffb1004dff89ffd50103ff94000d00230187ffa4ffb5fff6ff80004e00bd00610018;
    mem[647] = 512'h002bffbc0058ff930021002b0054ffebfffd0030ffe4ffb9fffd004b00340004fff0001e00080014ffdaffa8ffe2ffbbffee00670027ffbeffc300a4ffa70049;
    mem[648] = 512'h0086003cffa100f3ff73ff3e00d1ffa30089ffefffed00010076ff7bffc1007900050047ff57fff20067004dff6a0003ff9f00770031ff67ffcbfffeffdb0006;
    mem[649] = 512'hffc2ffd4ffd00045003a000affeb000f0009ffc2fff3ff12ffc300d6ff4affeaff87fffa003dffabffb7ffdf00af0002ffd70031ff400033ffe7ff65ff32ffac;
    mem[650] = 512'h00670037ffda0056ff89ffa3002d00530018001d00dc001500a100090052ffecff6fffd800350046003400e6ff4c003f0101001800790080ff8affb80064ffaf;
    mem[651] = 512'h00b10043002d00b600580036ffc9004d003e0098ffe50029ffef0029ffac0070ffc3005e0075ffe700b6ffc900330000ffefff5e00310005008800200043002c;
    mem[652] = 512'h000dffc5ffd3fefcffeaffd80043ffe3ffe1000d0015ffff0066003afff4001b003400470010009affb50064ffa9ffef009f00cdffa70097004eff9effb7ff75;
    mem[653] = 512'h004a00ceff84003dffa100f8ffd700beff78ff61ffce000aff8400430041ff28ff5a0099ffef0077004affc8ff9a004c0020ff9300fa00100011ffdb00a4ffe9;
    mem[654] = 512'hff9f004afff3ffc3ff650040ffa400310021ffcb003c0012fffaffab008effdc00670045ff88ff940080ffd2ff92000b00c2ffaeffc3ffb5fff30008ffb800e4;
    mem[655] = 512'hffed007d00050033ff83ff91007100ddff1f0068000a00a6ff90000cffebff5fff8b001f00950068ffc4005bffd900730095ff840020001f0072ffaafef6006f;
    mem[656] = 512'hff6dff9f000900e1ffff0065ffc00066ffd500270060ffd20032004a0035ff9900070011ff8f0078000fff99fff3ffb10046ffc30099001bff7a00e0ffa80034;
    mem[657] = 512'hff550052fffcffd5ffff002f00060054001dffeb004c001c0040ffbc007afffeff98fff6005f00530086ffa00002004dff9b0101ffcbffe7ff9f000affce00d3;
    mem[658] = 512'h0041003b00330046ffaeffeefff9fffe000d003b0040ff89ff9f002ffee9000dfffb0011fffffff4ffe20086ffc4003a001b007effdc006d007b004f0067001f;
    mem[659] = 512'hffac0069000f00a2ffcc0036ff4a007aff4900abfff1006b0008007cff7800590073ff9aff61ffc10071ff950019ffa8fff20073004a008c003a0072ff9400c8;
    mem[660] = 512'hffe30057ff2f006cff7bffde002affcbffc9ff8bff46006200900027fffc002cff65ff5eff72ffcf0050005c003cff62008e0000ffbd003d00ad0031ffebffb5;
    mem[661] = 512'h005afff0ffed004bff4e0038ff9bff90fffb00aeffbfff85002b002f0004005700060027ff99ff79ffd0002b010d0020ff8c007affc1ff92ff82002000200049;
    mem[662] = 512'h000f0009ffc5ffc0ffc2fff5ff5d00aeffe800840092ffd80085ffaa000000120020ffc600770043ff960047003b00640087005eff9affcd0061007fff700029;
    mem[663] = 512'hffc4000fff440057ff63ffadff860019ff82ffcbff91ff9200040083007fffcaffabff8cfff5005cffaa009f004bff770039004fffb5fff4ffd2ff42000fffee;
    mem[664] = 512'hffe2ffceffd9ffef0099ff62ffba002a00440038ffc8ff6f0046ffa40068ff81ffb900760069ffaeffaa0016008a0058002a000c005affceff650018ff22fff1;
    mem[665] = 512'h005100340013ffa1ffdb00b2004900250033ff78008affc1ff2f008d0039ffbcff83fff100500048ff8c006c002f0025fff9ffe1ffee006affc4001dffe9ffff;
    mem[666] = 512'h004fffeb00950041000bffd70014ffee0034ffcb0028ff9dfff2006f000200ba0015fec0ffe7ff0f0068ffe3ffe6ff8d002b0073002900d4ffbf002dfff9ffa5;
    mem[667] = 512'h00290009ffb7ffc7000dfff400990025000b004eff9affe300ab005d0079ffcfffed001dffbfff95008fffd3ff79ffd7ff8c004100cffff500deff9d0071ff9c;
    mem[668] = 512'hff7cffce00acff760012fff40019ffdb0026ff5a006c005affd8ffabffec0009ffb300010029fff70035ffd8ff6fff6800b8ffb4ff11ffa20032ffeaffe5ffc8;
    mem[669] = 512'h0064ffe50056006d0029ffcf005c005f0048ff560007fffbfffbff88fff3ffc000abffd20082ffb200220015ffdbffe5000f0083004a0019ffd00097ff950075;
    mem[670] = 512'h006d0027ffc400610030003cff800022001affd8fff10005ffdd00d70073ff620051ff2d000e00240056ffc800af0095005eff71ffa50061ff34ffddffc5ff4c;
    mem[671] = 512'h0065ff9bffc60022ffa2ff2b007bffedfef900ce0038001aff96ffe2007b0039007f0051000affc1005bff3affe1007bffe9001000380024ff75fedbffe900a0;
    mem[672] = 512'hff47ffe0fff30042003efff1ffa20043ff65ffdfff48ff77008aff8effda002000d4001fff7b002efff8ffe000640024002200d2ffb00040ffd2ffb7000effd9;
    mem[673] = 512'hffd6ffb80020ffae004900370058ffb1fffcff75002500b1000d009dff9e0036fff6ffbb001c0032006dffb9ff8c0030ffd4ffa900410020ff9fffb1fff1ffbf;
    mem[674] = 512'hfff8ff3eff620078004a0125ffa9ffeffef50160ffb2ff47ff80ffc4005fffd700cf0068007effc6ffb600110064fffa0011ff4b00b20005ffcb0024ffd7003a;
    mem[675] = 512'hffcdffb1ffc50028ffb4ffa10016001c004d002fffa4ff67fef2006dffdbffbbffab0009ff9cff81000affc0ffa2ffe1ffe100a8ff7a0040ff1500b2ffd60012;
    mem[676] = 512'h00eb0072004b00d50048001cffe3ffc1ffe60095001d002e0034004f001800a20041005100460084ffd20061003e0012ffb700f30009fff1ff09ffe20037ffcb;
    mem[677] = 512'h0094ffcf00ae00030013ffe6ffa8ffa90001005effc6ffd4006d00a3fffd0014006c00c60061ffd0007dff3b002900780003ff81004bffffffe9ff72007b0010;
    mem[678] = 512'hffe5ff61ff69007500fb001bff7a008100780094006000a20010ffa1ffcf0038ff01ff0dffcf00210029ffcd00420070000fffbbffb1ffda005300270051ffba;
    mem[679] = 512'h002dffe30018ffb20041002a0030ff900051ff08ff9a00acffdefffc000b00ebffb7ffb6ff7a00860052002effc100620077ffb00005ffb4003c0040002ffffa;
    mem[680] = 512'hffc6007b00520084ffcbffc200a6004affc5003e0076006aff9600d800250045ffc0000fffae000600110021ffe7fff600c9002cffb7ff79005a00130039ffe4;
    mem[681] = 512'hffddff9b0049008e0084ff99ffc1ffa8ffb8ffc10049ffff0077ffc9ff7300c9004affd7ff8200a2000d000700940099007500c9006b0003ffeaff4900070093;
    mem[682] = 512'hff77ffd40006ffdbff98ffc7ff9a0017ff89003d005000f5fff300590067005dffbe0048ff800012ffd8ff7cfff5ffc80014ffedff6affc800b5ff350001009e;
    mem[683] = 512'hff8000cc0086ff27002affe9ffa50088ffde0002ffed007e00ab0028fff1002d0090ff73ffeaff6ffed8ffc30038002aff83ff4c008dffc6008d0099004f0001;
    mem[684] = 512'hffa9ffd1ffc0ffbdff87ff70ffffffd3ff36ffc200a1ff6b00370080fff5008eff72ff8afff4ff9bffd4fff6ffe90081ffc0fff9ff73ffa4ffd5ffedffb00027;
    mem[685] = 512'hff2c0000ffc0ff240091002dffdc0059001100660039ff22ffaf0048fff30013ffd00069002bffb20091ffa2ff6fffe50034ff950049ff2f003bff9b0050006f;
    mem[686] = 512'hffe0002f0012ff5bff83ffb1003e0007ffed0008004fffc9ffe500de006d0035ffd20006ffc60056008d006e0006004d0080ffd5004aff6dffd8006affd5005d;
    mem[687] = 512'h0075000e0017ff7dffcc0071ffb6fff700240074ffbc0067005300b0fff5003c0059001500870033fff7ffb300860013ffe500070067ff9e0024ff81fff8ffd1;
    mem[688] = 512'hffc5ffc50014ffc5fff600090054ff9d0034005600ebff530025008d00270074ffc200900088005bfffe006c003f0030006a00cb005affe0ffbdfff5fff7ff9c;
    mem[689] = 512'h0037009f0048ff570024ffddffdefff9001bff89ff37ffbdff10ffc40020ffc20013fff5fff3ff9c004effcf003a006bffc5ff7affc2ffd60072001d0009ffee;
    mem[690] = 512'h0076ff2c0078ff5eff50fffc008fffd4ffebffd2fff300080053ff8c0004007c00a1ff93005e0094003900b90066000aff47009e000d003cff43002b00100098;
    mem[691] = 512'hff97ffefff6c005effb7ff470042ffdafff8fff20039ffdb00d1ffd90040ff71ff9bff8affd5ffff00160088ff6d00b60025ffec00420049ff98001f0044003f;
    mem[692] = 512'hffebffba004afff5ff7aff390079ffae005e0053008c004affc5ffb60016003a00a3fff10096ffecff750032ff890005004bff55ff73ff8fffd9ff98ff4700cd;
    mem[693] = 512'h0003ff940094008d003e0022ffbc0026ffe1ffeaff770094000effafffd6003bfffaffadffddfffafff20059fff0ffb0ffb1ffc8ffb9ff99ffdbff740078ffb2;
    mem[694] = 512'h0067002a0038ff84005200620077ffda000800970124ffa50008fff4fed80032ffcd0053ff87ffddff500065ffc000580068ffe1ffb8ffa5007affdfffbfffc9;
    mem[695] = 512'h0003ff150032ffd400300000000f0079ffe300ec00590077004fffb9ffe0ff21006f00630016fff1ff990008ffc3003bffdd0078005fff750038ff520000ffdc;
    mem[696] = 512'hffe7ff98ffe8007600490060fff1ffce004affc70075ffa5007cffb7ffff004effeeffd2fff8ff96ffe5ff53ffe9ffb0001b001fffd9ffd8ff3e000a0024ffd7;
    mem[697] = 512'h006a004b00cbff510067ff4900b1002e00330094ff93fffaffe5002efffcffcc00ab0002ffb900760047fffb001eff6f0072005c000dff4fffe1ff7d002dff80;
    mem[698] = 512'hff6cffe1001500a800250093005ffffe00d0ffd9ffe7006cff14ff7000190021ffdffff400310011008fff8b002900950010ff23006b006affee00650014ff4d;
    mem[699] = 512'hffd9000f004a00200016ff1effc6005e0001fffc0020009b0028ff8aff47ffe0000affd8ff9a0063ffbdff3dffa9ff450040ff37ff6fffe00034ffdeff81000b;
    mem[700] = 512'hff82ff5cfffa000fff8e007dffc5ffc8ff35ff4c001d0044002d005aff980079ff81ffd1ff670093ffddff25ff98fff0ffa7000affbefffe005bffd800480050;
    mem[701] = 512'hff85fff1ff9b003b002d00730064ff8b0000ff9dffeaffee0061ffdcff1b0015ffd5ff74ffb90045005700cbffcd0045006afff10050fff3fff70068ffd0ff4a;
    mem[702] = 512'hff370096ffb6ffbbffc4ffab0004ffe1ffc600430014ffb2ffcf0043ffd3ffc3ffddff67ff69004d0020ff860047ff7b00280022ff7a0089ffd3007effd0ff37;
    mem[703] = 512'h0057000fffd9ffdf0002fffe003cffa90011001f006e00250006ffd4ffd500290064009c00550005fff7ffe4ffe900b0ff78002c0000ffb0ffaaff81002bffe8;
    mem[704] = 512'hffbc003700260034ffeaff9f0028ff920020ffd2002a001dff9a00240040ff63ff8f00b10094ffa9ff66ffb50038ff40ffdcffdbffc0001400a6ffeeffb2000d;
    mem[705] = 512'hffe4ffea0027ff6aff7fff8bff83ffde00dbffe000dd00a2ffecffc7ffcdffdf00220043ff670088ff93ff280044ffef0054fff8fff9ffa9ffadffe8ffb30041;
    mem[706] = 512'h00c9005eff880008ffb1ff2affe5000c009efebe003000090123ffc5000effc2ff73ff72ffb4ff86ffe8ffb9007f0022ff77ffbe0016ffbd0014ffdf005cff8c;
    mem[707] = 512'hfffbffbaff900086002d0014ffa20078ff40ff610080ffbbffd000a5ffd40107ffa6ffc10059ff92ff96ffefffaaff9effe90058ff65ffc3007000cb0023ffdf;
    mem[708] = 512'h001b0005ffadffcaff79ff63002f002dffcaff2c00ba0059ff180048ffe40093ffef004bff6700040019ff740003ff8c00290079000d0007006d008e00300039;
    mem[709] = 512'hff73fff5002000040080005fffddffe3ffe90066009effee0059ff33007d0048005aff83ffbdfffeffee0004009000180058007800cb0032fff7001d0013ff13;
    mem[710] = 512'h003fffa6ff4b001f003b002aff99ff7eff8e013b0056ffaeffa1ffa1ffceffe5007c0044ffbf001effacff7f000100ceffb80041ffafff9b0017006afff4ffcc;
    mem[711] = 512'hff6efff20077ffa40009ffacff8b008600000025006b005cffc00025ff8cffdf0062003fffe3ff9bffad003400360030005affb700190040ff62ffb10017ffd5;
    mem[712] = 512'h005400200087ffb700880051fffcff46fff1ffc7ff8200db00390041ffb20078ffc7004b006ffff6ffb7001700cbffd8ffeaff62ffcbffba0072ffc2005c004b;
    mem[713] = 512'hffc3ffee000b004d0011ffdaff7bfffd00170022005300460043003e00270066ffb600000019ffe4ff9f00a4ff69ffc4002700090029ffc10003009400a6ff8b;
    mem[714] = 512'hffe9002fffb3007bffceff85fff700b5fff0fffd0095000f009c00e8006fffc0fff100b00043ff980015fffd006f00560012ff400092000b0062002e0024ffd3;
    mem[715] = 512'hffbf0026000affc90060003b0005000ffff40038fffb0097000d005300100060ffa8ffef0056fffdfff800cb00440061000b0054ffe7009e0090ffa100900091;
    mem[716] = 512'h0011ff94ff84ffe8009efef3fff4fffd00abffee00540008ffca0064ffd7ff95ffb2ffebffefff83003a005dffdefff8ffef00720005ffd7ff4b0005ff9affd8;
    mem[717] = 512'hffe8001dff2f009800660035005a0056fff4ffcd008a0055ff87006c0045ffddff3fffce0041ffc10025ff8cfffd003a0063ffb8000effc2008600efffc4ffcf;
    mem[718] = 512'h0004fff6ff8f00310033ffbeff2c0038ffb00036ffea006bffcf002bff6900a3006affa6ffa600810049ff760016001bff9900c1ffc4ffda003e0030fff8000c;
    mem[719] = 512'h00a50065ff9bffa1ffd300850030ffb8ff59001100250006ffe10057ffcc0016ff93ff7a001e003efffe004b0012001f00ec0038ffbd0041005e0005ff3c0033;
    mem[720] = 512'h00980003ffc6ffd30029ffce0041ffcafff7ff8000a4000a0043006d0059004000220098004eff8cff36007effe60029ffd70003ffb3002cffaa001100620024;
    mem[721] = 512'h00a20064ff8500370037ffb400900089ffe800d60021006c001800900052ffd7005800a8ff3000780020001f0014ffb70044ff70fec3ffecffe5fffc008900b1;
    mem[722] = 512'h00ab004300240007fff7001affdb003aff7effeaffb7ff9e0006ffdc000100000022ff840060ff52fff70087001fff9d007b0027ffb5009cffcc000b0021003b;
    mem[723] = 512'hff2c000affdffff20057001bffd5ffcf0015ffa2ff25002effd2001200340009ffc2005effccffb0ffc40020ffd5ff890001002eff9c006bffdc0054fff20055;
    mem[724] = 512'hffedffefff4800a400250026000b004bff5fffd0ff8dff0800b9001f0035ff83ffca006b003e00e4ffd1005c00b1ff6cffc4001700aaffa10032ffedffccffdf;
    mem[725] = 512'hfff4ffe0ffa00002ffc80026002e00720068ffa8ffe1ff8b00380050ff6c0146ff97008dff800024ff64fff4fff9005eff6c0019fff8ffe20004ff92002affd1;
    mem[726] = 512'h000cffdaffdcffe7ff6800ee0028ffcd008fff7dffee0044ff75ffe1ff550081ff75ff71ffb40029004dff32ffcc00e2009700a40052ffed0046ff8d00010077;
    mem[727] = 512'hffef000d00590073ffccffda00560069ff63ffc7003300370014ffa1001cffe7007c004a00720014ffdeff860054ffdbfff60031ff620025007600a100d7ff49;
    mem[728] = 512'h0070ffaf002bffb6009c006500f20034fffaffa4ffac0077ffc0006cffd7ffc30013ffd10005ffc1ffa6004d0091ff91fffc0012007fffc8ff9d00beffd20004;
    mem[729] = 512'h004c000f0055ffcfffdb00acffb300750044005bffb3ffb50004ff9cffc1ffb4ff5fffb6004aff60ffa0fff8ffdcff5e008fff47ffd1002bff8f00200011ff94;
    mem[730] = 512'hff880086ff79ffde00280108ffe7ff5e012d0068ffdfffb500b4ffef008ffff5ff870098003eff940043ffddffdefffd00a5002500320050ffe2ffe5ffea0021;
    mem[731] = 512'h0109ffc70052006effecffcaff89008d005fffb40078fffb00380080ff94002100870036ff74ff71ff23ff50008100380073ffec00540054ff7600830059ffbe;
    mem[732] = 512'h00a0ffe20082ffdd00210062ffc300520039ffba0063006c003effc3ffce009cffe6ff5bfff60063fffd007a003fffdb005e0057001affca002bffce0073001d;
    mem[733] = 512'h004e0021ff8ffff600bc0040ff7cffdcff6f00d4ffc0006e003bffeeff56009dffbd0019ffd7000bff91ffe2fff7004eff8dff85ff9fffa10000ff51ffb00001;
    mem[734] = 512'h005c0014ffd400cc0039ff5effbcffda001bff91004d002000520062fffc00af005000630020ff97000b0055fff8000effd9fff0001300a200a9008f0042ffd6;
    mem[735] = 512'hffe90086003c0009009100d9ffa2fff1ff8effd3ff50005e007aff7affe90050004d0031008fffbc00f7ffdafff70021000800580021fff400510027ff69ffb0;
    mem[736] = 512'h0001ffd6fffcff73fffdffe4002f0046005e00a1ffccffce0018ffacffd70088006effcd0035ffd50096ffc10023ff890060ffc10071005cffbbfffe006b004d;
    mem[737] = 512'hffb2ffafff450044003affacff34006e0040ff7bffb3fff9006dffd6ff58000a00320084ff7900a9ff9c006800520017fffbffa9006aff82ffc9ffa100090022;
    mem[738] = 512'h004effa400010051002bff3bff74ff340003004cff8b0017001d002bffe1ff9affef00180029003fffc70049fff9ff8fffe8009f00140031ff1f0036ff64ffb3;
    mem[739] = 512'hff910023ffdeff280058ffbf0087ff47ffd9ffa60054006100190032ffaafff3ffe70010ffd2005aff82008e0034ff83fffb002d0065ffd40071ffc10013002f;
    mem[740] = 512'hff5cff6a00120030001100250028ff91003e0044fff9ffbc002dffd500760037ffa4ffcb0039ff8cfff4000f00770075ffbcfff0ffbe00680020ffd2ffc3ffea;
    mem[741] = 512'hffee00940029ff94006e0094ffe80097005d0062000b0076004a007dff7fff95ffbb00b8ff3effca004d0065001b0048ff69ff71ffcaffcdfffa0073ffcdff7a;
    mem[742] = 512'hffa4fff90012001c00270090ffbe007cff8a00eb008cfff1ffb4ffceffb3003d0014ff4aff35ffa1ffbfffd900100078000d006bffc2ff8affadff3affe0ffb6;
    mem[743] = 512'hff190029ffefffd3ffd0009800350078ff270012fff4ff8dffab00a6004b0006fff7ffa90021ff9d004200360022fff2ffeaffe0002cff4c00650029003bff28;
    mem[744] = 512'h0076fff3007cffc50060ffc3006cff87ff510094ffce004bff78000fffc80067ff95ffeb0092007e00d70006ffc2014dff540009ffcbff6dffaf008f0051ffcb;
    mem[745] = 512'h00b5ffb2ffcbfff8ffef00670047ff910041ffd7ffd50025ff63ff80015efff00089ff8f008cffc6ff8300af00a6ff7fff73fef9002d00190041ffacffdaffa4;
    mem[746] = 512'hffae0015ffa5ff7eff89001c0013ff5bffb70087ffff00170022ffc0fff4008c0001001dff810009003fffc5005fffc30022007c000e003fffae001eff96ffb3;
    mem[747] = 512'hff99004d0040ff4f008fffb1fff90013004c008700de000f0052ff7c002e0003ff9effc500a40049ffbdffc9ffe2ffad00160025fff4ffc6ff9c00000075005d;
    mem[748] = 512'h006e002e000500de00860053008fffb1003eff0dff5b004dff79006c0069ffcc00dbff7fffceff9aff58000000240006ffb3ffd9ffccff460038ffbc00330077;
    mem[749] = 512'h0071004fffcf0012ffdcffc70036ffecffecff80ff9d00200067000c0025ffd3ffdb00e90085ff8f0088ff82ff87ffd400000011ff8f0019ffe8ffd70104ffea;
    mem[750] = 512'hff6c00fbff5e00b9ffb5ff5eff59ff37004700780014ffb8ffdeffeeff7000b9008900710000ff9300540019fff9004f004fffbdff520064fff2ff3c000c00d6;
    mem[751] = 512'hffa60034002bff83fff9001d001aff97ff76005c0085ffeaff6fff13005cffef0133fffeffa0ffd40078ffb30036ff81ffacffa0004b00b20042ffcaffbf0015;
    mem[752] = 512'hfe9e011cff93ff36ffcffffbffba001d0021ff13005b0082002fff9300f00042ffb0ffd9ff57ffc5ffd00003ffd6ffdc00ebff430064002fff9a005affcbff8e;
    mem[753] = 512'hffcaff94ffa0001dffaefff1ffbb0016ffa3ffaf001cffe7ffb1005dffb9001200570065ffd400b70090ffff0074007f000a0081002dffa00024ffe7ff370057;
    mem[754] = 512'h0008fff0003600110034ff4500160020ff2aff4500ce00340046ff9c00430044ff51fff100530035ffc8000e002affc20026002300efff78006a008fffe6001f;
    mem[755] = 512'hffdf0018004efff8ffdc005c003200b6005bffa8004c000affc3ff34007bff910013001d006effc2ffb7ff5fffda000f005300e9001d0060002a00a600600045;
    mem[756] = 512'h009c00640006ff72ff840020ffea000fff6100edfffa0037ffccffaf00710034008f007cffbaffd8000c0009ff9eff7bffa6ff640029007500660066ffc70076;
    mem[757] = 512'hffb20049001a003d008500430093ffe6ff9a0028ffb20054ffebffe2ff7cffd10012ffb1fff40058004c0039ffbdff6fff590018fed2fff2ffc3ffd800440026;
    mem[758] = 512'hffbe0053ffc8ffc6fff20067ffd50091ffc1fff70003ff90ffa6ff9bffe60077ffe3ffa40003ff65ffa7003d0053ff85ff81ffa70042ffc0005fffd7ffb700a9;
    mem[759] = 512'hff64ffcaff4affe0000bffdf0011009dff7afff3ffdf0048ffa5005eff73ffe2ffdaffcaffd7ffe2ff93ffc000dd005c0041005c00b000a0ffe5ffe6ffd200c8;
    mem[760] = 512'h00300040002c001dffcdffcaff32ffe6ffe7ffa400510002002cfff000a500410037005b005eff90ffd0ff63ffb6000dff82ff2a0078ffdf0094ffc20001ffe1;
    mem[761] = 512'hff02007a00d000c0000c0001ffbefffcffcfffe1ff7f0085002cffb700b00077fff4008e004d000ffffb003bffe300ee0086ffbeff79ffccffa80088ff71ffd9;
    mem[762] = 512'hffa0ffaa001000380029008600bb00410012ffe4ffac0013ff880047ff690024ffa70034006dffc000d200ca002500860043ffc3ffafffcc000bff68009c000b;
    mem[763] = 512'hff890061ffaeffc0002eff8affb90035fff0001d00120027002affad0017fffe007effb400b2005fffdeffe5ff9cffe1ffd5ff9a0026ffe3ff51ffcdffbe0086;
    mem[764] = 512'h0054ffb4fff1ffb7ff0aff07ffb10009003b002affdfffbf004effcd00b900260043ffcfff9bff05ffbcffd7ff870086ff3dff3ffff6ff9efff10047004b002a;
    mem[765] = 512'h0037ffc4ffa4ffaf00300005002c0005006800340038ff7cffa2ff6300a60081ffab00910042005e0067fff8fee9ffb4ffb700da007a004bff4300cb002d001c;
    mem[766] = 512'hff51ff55ff92ffe1004dfffbfff4ffc10029ff6effa5fffcffcb000a004a000cffc3fff200c8ffdf00360027fedaffaa001d0043fff000d0006100100032ffce;
    mem[767] = 512'hffa5ff78ffa1ffb1004500050016ffd6001900c0ff980000003c007f006e008c00adff98ff900037ffcbff3effb4009700050031ffd5ffdf002200720078ffba;
    mem[768] = 512'hffef001c0006ffa3ffdd00700031ffc9ffd2009effe30065ffcbfff8ff8eff92ff760061001b00620075002c006d00400022ffe6001d003a0032ff6b00a5ffa8;
    mem[769] = 512'hff55ffb2fff20062004b0019fea7ffa2ff38ffdb00c6002f00230081009bffe2ff85ffafff40ffe8ff5e002e007d0074001dffe9fff4005dffabfffd0011ff3d;
    mem[770] = 512'hffe4ffd1003c0037001aff7600090065ff9c004600690094fffbffcdffe60034007800c4ffe0000effa0ff23006b00230075ff29ffa3ffdcff8e002b0053fff1;
    mem[771] = 512'h0094fee2004cff93ff8efffffffbff980030ff6cffb300890094009a0073003bff770015fff90055ffabffca008dfff6ffbb0040ffdc0001ffd7009d0065ffcd;
    mem[772] = 512'hff540006ff6b0063ffab005eff42ffba00a60091ff72fff10093004dffc90067ffffff91ff98ff4affe3ff84ffa6fffbffc6ffafffd70036fff8ff3b0033fffb;
    mem[773] = 512'hffef0042ff9800bcffe6ffe600cbffbd0022ffb9ffdd0027ff78ff60ffd0ff56fffaffdefeed0050ff9bff5fffedffdfff8afff10007006f002600830055fecb;
    mem[774] = 512'h001a0037ffe4ffc7000400630019004a00440037ffbc001b000afff6ffdd006c00330070fff1ff7f000effafff8cffdeffd5ffe30120ffeeff95ffe1ffde0030;
    mem[775] = 512'hffc8ffe9ffdd00530053ff600048fffdfff3ff97ffd2007c000affbbffa5fff0004e006d0011fffeff98ff5200340082ff4b0061ffc90029fff90049ffa10035;
    mem[776] = 512'h0042fff5ffedff06001000b7ff54ff73ff7cffe1ff9d003cffa6ffcb00590016ff7dff3cff2f00610055009d0035ffa1ff9b007bfffd0006005d00470043ff65;
    mem[777] = 512'hffa70090ffbc007affa4ff8f0009004dfff8ff7800130039ffa2007c00540026ff8fff78ffb0000f00a20028fffd0001002b0059004100b0002a0012ff41fff3;
    mem[778] = 512'hffda002a001d001cff62ff5e00500064ff9cffb4fff2001f010c003900b1ffe000cdffac001e00a0ffdc00bd002100190039ff84ff140054ffb6ffcc0000ffb8;
    mem[779] = 512'hffd000bdff77ffd8ff71ffdffff1001a0008006800370117ff8bff790038006dffb8001c00120021ffdf00070042ffeb007500c40026003dfffc00160091ffc2;
    mem[780] = 512'hff85000f000fff60ffecffebff65007affd0ffe0ffb60026fff9005d001cffb6005d0098ffce003f000d001fffc9003b003effe7ffc7fff3ff430013ffdeff63;
    mem[781] = 512'h009eff87ffd2007800340069002800d2003bfffa0090ff83ff7fff7cffffffec005bffd2ffb40058ffd1ff4100010016fee4001cffd8ff7fffa8ffa20005ff5d;
    mem[782] = 512'hfff9004400610080007c0054007dffd800b1ff350090ff9a00250024ffe8005aff4f00700020ffffffbb001a006b0016ffd9004d0006ffe8ffd6ff9bffb1ffb1;
    mem[783] = 512'hff7400ca00020002ffe90037000cff58ffd4009800a60051001d0036006affedffc7ff22ffbfffbe0097ffdfffe6ffe8ff82fffcfffaff9b0003ffcf006fffcd;
end

always @(posedge clk) begin
    data <= mem[addr];
end

endmodule
